`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
p5MldIvdMIoYJJgWrB/HMO/6Mueft2nWeMyKdzdicWmOMpKHpc7SwddK8KXaTOyj
ZrVtZuM2v6HvGAC77mek7DVPhC5Q6LhQdhrKbs8ffsUaWhWunWgWSHE+sSdUOV4L
i24CSrNUUtJ7o8sGPi4Q3r9Xeu59fq+qkVlLaLTrOqQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3264)
5YTag39o8F++oP6rpOVdKbb3PwcCELnv3L5K/pO6wfTzbYQ+5gCya8AlyN0tLVAJ
g8W8eHPaslOwMiXUP5a3ov0JjFlpa40FjnVyDv5DkbflZH8fcK3Ng7o/LY4g+CQQ
6GGz7b35UkuW5PScmXbuO1EcsQEleELbX9x5xJNLHKxRwZSL9I2wAKxMIxGPxlel
Q1NO24XOkuEwnsG+QPqcPneMy84sLuFkLHPeRal2rNLPeR4IfEP35bSIhJZmJOik
Drcypvs+VDZy5uSaDzuQA89V47ARxkTRaMDa5kFX+jFCt6RTc4tEiMHWxUnt0RuS
7T+zmQUCR/ybikXb6t6zDDuUmS3EWNFT6+oL5xXW35WDHyVo7kFRJpwf6lEaiDP6
vqErBzHwzEMWwdr1d/BKUz6NNMvYaMQCJVg383JFMFC38hH7AL6EJEJLaVVYu828
vqvoeZ9pXtCOJLeLJNHNvkKFSUP/6E7FKvSU2iHTbUjkKqm90LEpBUCjH+kIpaM/
yL8Yu5gXHBogOai4mMkKSxTCxCz1X8VCWS5cQZu1+z83UAzoKaljU0yJatLLdTyT
8QTc436Fj/J8y3Iwb161Z67HjtSa1tsg+w1quLfgvpY2sncO0X7FA6DNTY1JjLCm
AGMJNMBRqYZev1ksVfME+6tnlR/ixXcYYNoXpPwIaJIDgsARhsNiRnr4IUs49FKT
HRkhNIbxcrGEGftiLNHZJmb+x9oHXf578Thoqo65YYR6bXS2c8qrAkkdysJ5jfoe
Dgwrej3bb5sRtHTa4SnrVSEjVG6MMwNWmtCL18CciXZ7d7+B4Hxj0uXGu+9lX+3C
+JWxPaq9IuRolYgLyGpcffAd1aqRC7BsmQ8sMgV4HqP/rOD/GXb/t0PWJwfcEqBq
okvNuD/f9vej3WaIk0I1mSE3yxnZZS7s5lFRtScH9cywyROTlXoMnBugdOmUwpVd
CpjH5ao03pXgpBB1RmuIBWOV67gUhgYNTKfxcnsZOdZ1w4VpgJOIw8eFkKVF2Blj
TgRr6IBMhpHGNms+nBdRpFdJ6sdtCoiE+GEyxdUWc2jANui636mt6HilYVJ2chFd
v/DtzwjEhjN6TzaWct/ikJErSdgAIpC2NYynGcGishwwC3I31FfssYB4VG44G6zz
SFjUdXJptOMNvJZDV5Riff53snBzx48qLJMJjVvVu0dZ+7pVbwik/JpdZ53QIfe7
TarpMFkhya4o7c0CN85ic6hlhz0cMFFYiBLD1ZVWeoNsYOj2SLhJNAXpPajEMVF4
C7/XyGMFumRyna5MYDdpO2cpmrEQyW2VP+87G+6x3yN3KaqSIPQF6C5NjT7gJRsY
R4kuIluyyU6qyYtLVGTNUySpa5baPKWAoi6duPWHWiODV68Wuo0UxO5SlAFYTYHj
rOHMtGZmGGBVC1dB1JZ1/eCArSX0aRj6aiXI4FfTx8G6Sxy3H8rAk+gcItr7jjsM
Xl8ROZHUGjwh3GfTCIRZFaiJweaawEM07N1XunlmiX46AeQYFdUkzAonOpHlpT3X
NurhqaWxV8W5iiSsFH/5hGptqvW4Qr7IliKfsDdKC75OH5Q14ifgFWytHJhJvw5w
SBcoi0WcH0CWyeyqK0O12JFwdmTa+j4MbCKuFYA2JmveXk2ouZpJh8SADJZFJXIV
/mQ43iZxxcq2V5/4zUWhT0+02bUjgceFeGYR5mNA3ifWs1fwNdyKieLpJhyQDZHb
qZbmVlBy9AGO0bqUUvZODzONuQ2hz0SodhBwAvLGDjjPCkMIV8rLskQUGw3fj2Ru
g2lYAoXX3KCdQonpUISSUFz3P/O4yffqHiV0Z+OLa6uFdvoXCYr/YBlXyVZIffB1
e9XjyKOTbcHI5Bx8Dcc138xRwJlWd7i6KTduBtx/+E/qsgDEWZTcMtEms9vPuktc
y0qim5lmp//qu+Q1eK4gAGCh1ZhTx4BfIpdFNCUQvF0HdShXj8Rze0zsDwtWYULh
mywwveWyUkOeXXDkskU+V6kKKObqaJoTabJh/uBpjIzYoy6FDzNaVRd+uwChQrhH
sKeFkI7ccdo9rbvXdxJvMKSiR6FJMfHU/njOm58QhUM/E6Pf9a6XMgq/dKj7HsA6
wVyYgZyp4mobAK4/QyDkqHnnMHKm4nS2sKregvvuOwuT+xXStuRSQxbcAEuUbEs+
fVulvvBGkFodwePaP3+wT2VZiA0CJdzBmn00fzxCctZ47fDYayesQpNltTeolJ6D
ZsI8JAE7SXYimSINRn4zmw+/pLOa0gffPQzMryVaLf/4Oz/O9P+/0fDd2mwap07f
zENm6TxxjP5xnCdbWNa7wuuYd+n3nZdf2C/ELUeeuBYw7BBHLoebE7jXcT9FBmmV
WAPnoCqdcexaYF+BTmMx0eNW4vtINA5NfqXOhELmy5agOYnucBHKCDlWrkz+RNjV
aXaumx15iLQz5JXebesZEfI83DOqPybGGgQNll0Dl5i0nr6s1DhwGi77uiYuAS/Z
7lSNXix/n4aiQ0ninnRkc9jQL9pM5LQ8ytZqSfxjOLCePRs50Sorh7G2J6JbX4iN
ImuFgjESv4k5UQBbSnnoKIsd3IGhXOzfsWZIQTCKx5c+jUyG7oUpF8havB9WbVq5
hyHFxgtcL/F87PCFY9urb5Bl/E/yWyE+XjJxSmUATs5LMOgM9H0G+sr9ThmBNTmB
DUCOhOVKI/FJwVDo7QV47zCf5v3ho4NDWCh8FAUXASc+cRhDUVw835SQf+0iPQrZ
dITnvZGgRepDdVChcgbu44iZFVwJZSv95dcioNqPP4jH05TEOCbivuI2GplWm8Qz
FSyr5LNx76Q5/drLwPHZcCpF2FglwROqqVX1tBHPNtyrqzpQC/Z0V+8tCV2SAte0
IISsUwhSDdTyqigNT8GJQuzPavcPMBext45RxWzif98P8GyheOAvbWeuf4E3vP2B
r2gM5dveFjG89JMlO2rCjEGCIgC/LyWkkzhshdm7kpLAy+s83jqTBQVt6fkvD+jq
arLgeG7uT26nnNxNxGbkeJcJlYBadCaY5F8TmhII/nB3/L2NmDMYfc+BoWtVbVqp
kzMY+WNQYWoAVuQ8OQcwoS4A/08Ero/RH8F/bTGmzOGHgld7BiZXAEJjWku8x66u
mhNrIRqkj2e6eGTRhz7bNIrhAqy4bSbWfVJnZJ4+KeJXXqoK7PcUPJ3qzaimJYFf
fMKMNSbFZwJbgv8BfkC4/y7qdydmZfPqnCTvp7gxQkwVe5PnFxlpEVvM95gYX6lr
fA39zmdvkb2RL3NEvh3PATXgC/4UONsr/IHGN5841ZXwk7aAdXleuuJoVKIQP9Al
J5q1+Sq26vo6+wDv7KYe4l1OnJrn6qqiynkEeCdtnMOn+jxp2Dgs8GWDEJhnl9H/
j0ximPR3qViF3flfsuGYSDCc72+3y18Mj+mFbLI25N5T5Kf3A/BSgIiyowvL3JiC
36HKxqHKMuGkg/+txUSQQc0DIYuAlMH9Qzr2XEZlUA+N+NrQwLvrARYmKMMfx67C
CtqKCuNeKy4c8enE1RjNaQjHfKCbqeMlNyzCspfTOGHOomyiErc/5vDoPp6GHEt3
766hUpVrgVvhuCFYt+YZhQ52Vnv+gZbwTrTReAtNynj5IMFdiM74Jx+1XAfTP145
8CzF35jMZkMxan2sJR3V/MUMR7Dryz6oS/h4/4XZ6ZDukKieKzDQrqV8yY/77I4W
04yHYb5xEW9dKd1eRyb1NY716uZJboNkPemPPTkrYnqE2IqJrsX5u/KH4itgsOaO
yeE9c9GixVYfu98pDL55Zjn9p6INZrGFAFZqrgEC9eWnCzo16m89KjNMGjt6h/qI
RoUKtqV96fBfKi9FSLUKXDHrJZMKN1GagEdBhKZjt4WWS1ZneuYutyvtSKv4RZz9
kNJvf28o8HKPr8FZ6Fe8beWUa6a2i62L7ICqFXZN1ITyQHKYnNZ7r40GQGXnRjI8
Sjhu3dThl3a/w3wJrvbETidSiY1Mmp6dOXq9rC25eWrRvmPZghqBAczR2J1/nf4b
sfkZegBALVkH12qTNzj9Sgr3N2dhP/Ykdq2YX2OwN5kc9+VDA4WTwW1okZjmtojV
fOJ2UTus3mv1jR2avSWyDf6QboHpn44WwHMigv4m0ZeGDlyDJmMA3JkTHWk7unGB
+ZveCessVqd10LRDVI8ffEsZryHP/OTP6i9X5xbkOMyGNQZlf8D832eOcBbwo6Y9
9O8VgDh9LUrxjrZC5HNLOsRoFgvqKcFdg3bUmxCNu5Y4Fk8TPEMBgpbePUfkH1jt
fpyIMniThaul/ZaZdBmaPZ0B4cw0Jde9Cz7QzQkcOSOaIcJbd0GstybKTz6lJYce
`pragma protect end_protected
