`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
by55eB4XyP7wqUHY66LAjVZ6WpfTTRHxpFOmS0GW2m8k0D3M4wuBU4yBquNQAy4A
64z6Wyw6jo2SunV4LogaG4R6Ej15aCgUBOHYYMW+zcIHOo6cFGzhXvL62gMU4VWS
FgqKEuFFHFfNDIb+AN1tTzhdCpjoGEUY2plH4xAGuqg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5216)
Em9G0Bq12FjWZ5xDV1Fxb5o3vHjJBzvuEyEKzx6gh8f2BX1Y52Kh92hysBAC2nab
5K7WzF3xU2iopNFpgOyVOWtDM/xwtjM5xS/ZqlgS7sYudoeFt5qFnAijTjb2xAj9
IqhenhYe/dE8VnjWtzLyZbFnXYbnbIywLzAT/3h8pvg55ven1swN/F7CidT46oDU
eyH2lvs/7LpGdQhM906CHQF/lNI83hqxeeWii6PJncNH5UAl6aZ/4KAWM2mYyn5C
aXtTFAfHXo4+J/RDDQpCWY+B4ZkxHuEamkzs/S56db//HXfZBIiPDVrVIF4IFcYB
JTcbdDcdO0TXWqdUb5Y3IJlmr721ZCkEJfBC0II0QeRxyzUK6QT0jp6a92G1PoDQ
qKbKIRrKq51rqz7G6LwPtVjBWNug/fW6TirtYUyVsMVV9hik+YSblHWzLylTJYWf
UIxr+pT2k+X+10PcolMLzHdcuQc4FeB++8c2mN3/IJ3UbRH/E7VwswqU0kIoKUTe
IEEksUwvt+1AGrbPm04iG8u29G0khPlOfE/0wlQfU5BiuwSrspqqym7Q39bdwkAr
7vKXB0DnZdp7yvlnNAsTtozohH2+F8A3tBir6AGI0/Gi5kU0xDEAaqa+XM457KGI
+APkgyioqElQyXr4xRc/uQPqEPR1OJPoGZJ4XFQdib2TpUrY3c+zxtVv7c0h/btl
9/M2XBCr2jJLNLQl7MGEncQiFKTv8ePg7zRJHOMxHJbrVpL9YVmcBqoatC6zX8/I
EX65QY5EB17RprjuURNDeT6lssKpriUp5drC/vVAjAc6IpsgWTXmAtKAhTP5qrlA
Wc7Xw5zJRpAIX2QIW181AODgs8yU0SaHOr2AyBiHeKyExFIRV+EvlXyJxyUF0vfN
ZoegwwxIV8jPHlr2JWicViPymGJddH5eBNK8BFiUK5+qz36N4TtsQQbCw6Sf7d44
BA3P3yXULj2fXZHi0r0HQHlxAZrcvN5JW2oZ5QLy1dX5JQMHhzY4ZwR6L4VZU1GA
krkJ88ZLno25mkS96/f1g7nmteV9krKXW8vQETQeonWv6O7pAPgpgWp6sSGK5i7u
5S36vHEVV/oVnMkjKqM/q/IbNNIpXR7BferQPl8JzRQJ6xAruYxdyGdKGixwmOff
jkQ5m/56CHEfOGEIpVhzDJXF2tck/ijL+d2P76pgx8RboPk3T+EV/KAH3zkZGhmI
2SxKDna36n73+0nAUxFJHHaECZ5maX6uFmOp059r8th0zJFYM8mMFhNzJQVRoBsR
n04qwPYaf6uKfdLLVCUUQZTNgo1epbv8Z0muUJe1WB4tdSAYLRsN1aS0/VfYPFdq
qMSQe8xzBfVp29mu3tOGLmQpvxstUtSmIVipPpvbUvgGSJpRALMIMMqUpCoKv6tB
jsILCp9LCmM+3LXmQ3/UhcRRgZ+b+yILMEaFABsSd0YuESq79u7/7raWI9RXfkeK
0+7+ozZhz7KnA0vk8yTarvWqSzaxqrMDlxazAifJGEpudGQw5H5pa9poyT3RB0gp
zw+d/z3gVLxEln3/ojOAgm8gaPkk4upaZXF/S3/bih+GMmZcwklCUmCbbSgBioNG
l2ZdK0ZgOdaHJKtDrYlPCctAByvP5x0M+lbgbCYpDzm+4Llt2zmSM9eVY08sJQje
aRlRKROgJ4Yb0Frl8WOYMhJ/iGMcxJmNBGUbJR2iqr/6bHt5Oc/FYSONcjYI2CjA
4yXpZfh3taO8oS9P6fLfvBUtSx3Rv+V++f8U+guN0Q9yjsNiy+LSghjpuB3ki0Gg
93UC7U8JK0sak1MbuK0fmYv42t2MRUBCBN5ce8AgxmxV8urDBBVAKMh1j/X8UDfM
A1dLD3Y61SKdv47nAfwupBybUhqZvnkA+Kd6jMGNeK1Sec/d4KkEvMqTyYHxtC/k
7DQZLCp+vCnn66Oj01rtP2VfPLvSCTJKWA/WDAzR80jfzgnrUsCYAxYKUTUKcPkz
zRt2LxaTzpFVyRygIFQji01zbE2HRfTVSBGrR6OKf5pKOXAy05WO1AQAiV2xBJPI
mZFBD4sSwTBTRj4pYgF0GcVMdfC0s83rmPxRDyRtsv7JWHU6v0vcJJCU1ux3zWUa
qowG48gWuboYYsoLKS72NTa2UZEboKy1O28hMC7Gzh83nY1iGXVbgbtuYPDz2qFJ
SAqy/Uw2sczR3+qxZlFk5vX6iY/peVT4JzjUb8wT/Vqd0ZLADmC8d5sQXV3LU7dt
OwXioebHcvOIJnkHcrNS32bhtHFkkGspiv/YPXHPAeXPzfVoAv9d+rjByMd66sfn
p5FYg3ySMZ0NXFmm7qXCTd/SZ90zx8clKwjh/wzTrUaZ+jEyPZZEebjyKnORfTCo
MJCp5LW7SRDK4KltLBRjKGW6/0974wllCf2zueeo8S2Zz2h1FTRcm8XLaeIJA6Y3
ImO/0BpuXy0LOomuUEEtdn2F4ercNK76567yDW10wcKfc49KhC6UYMFMv6P5TMBO
tloGsXX3dEbWCabKtwjgQSNBJV2iRAM/KrKk9qu2QEmhLdFiM7cEZc9SiqfPMH1h
RJUqF1LLx7zo7Nf6EY3Cwc3p6XPg3oy8U4LWvbr4K/68gDZJMmRhWuC9Xx8W3CMr
9B/Xq4/wYQUZ/KnncyUjpMxVx257gsy13HLt/UY3q248XX2zaA1+lirNGuIhz2c+
9epC3onq5KyvcGX17jClzk8QN6ExIy/c4d76oBLogWEi+fujuXP8JemhwOyvlVvL
sKXD/Sriv3+D+I0hQuQJUfseiUMKRY7cMCXa/GFMg/w2gVweJk4MgC7kJOPAcGSB
orWqtFPWIDzi61JFFuahi8JDY/KBB9FttDIHCFIDG+n8crg0IPrYkv28C30BBOsK
HooXUvhyw3dztsF2m2bmlGwEvat5cEDdtdlisJmzZuP4Baj76ug4Db1ErY18n55h
olhLc9LRbfuv+Y/z6+ByEN/JviHWYwnHkJR1xdRQ2g+za8ndgBNbNdWhNNt0/IwG
FQ3XXTo+rGTCMdlc3kfPYJnCAJpHpQzF7cl1dWcUEp1ljupIJ99bPo3ukJQkfx8x
gtgkpyNB1eml1nB9dF0nqxC4RF8ZF6G2J0fpb5eqiSS+CqAOfKA6V7QRDuFr+hei
qoe9jM5i1LXi60sg4rLSbVzjhJ3Jw9c3mWzlR0voifFaZVAKsk5GiGG9cv0YlgaS
alPfD/TbJMoYlcWo4mYOF80xRBf0Cu7P0qfGqXjWqR/qgDNZtGBRhkoZ3FRYMRnn
q0Oo/sHzig5gr+qJ0V/QgVgh8BN/UN0vYbvNR0WhcDIh2fbSTWCrnUM4lBVbZucg
j5uIHpS+mz9gboTUttOeKzn/sv3sc/wpoPGSp8XARofeWukGf1GCGEnHXqSwS4hj
pQlAt6QhGkv4yHkCq/6RMbS+l+hK5ZyZDLIJoKB2F2OiWJ0XM31wRvd9w32LwAbO
yc5JGtBdre/utYUBH4Hq5uXXHJmzOkBXG7Ts3L8N4BClAU28I9idLUm0yZ4dR/DE
hk3CevefjS4NJnAjANHIZqdQwRIurFqyIrrMgyVOL/OrodvRnP3iBrUTF7oqi++J
+kvTe+0qsKa1CMCswZHnXkiJjml0ILJORBfeR0R8r+zgmc/67td5itdB1nzgi/Ny
Yy9+2BfQczXtalGir8xMcQlsI4i+PhFEv870pBd8EZdN0r6jPTuEG1AqclgTjHOK
vBMg5c3w5AvtvQAFNzc/YFEfw5dKevUi+6WMRo1anOeXY+gp4Jm3QBNw4vtxhIEK
hJjptpGcacqrjxgzO7jOUuDzZnwuDjOs/kGbx6w+sCjEcSjLjrWD85LKR8KJaRpM
p7gzt3cyuXVMuE9GW40kIqpmZLqEmp+bDLMw4CIoesc3WRypCwV3rxXoTe6jgloX
pby0pr9/PGd1B4fYx8P4N0IqqOgR5qRVa69EQKQzTksuPkl/gnrRgVf0tXaw4Ptd
HNVJJUKgxUHDuQLgU0V4eeJIC+YbS1d6UFwVljqSWghF7X0+vtWUiUOMuUULDr4V
Yf1id6iXnO1pTzPj51qZjgc0dhYoeQZarThPmZSxGM512E6sqSAhovQOcLgsWYPM
RNNUrNPzxn/XXXaQRWMf0RivX+QCUYZLUKX3p+5dv0ca5DquKzjrHCShr5fySwrD
/x17wontG38ZB6EPDC4mjf/OBUPPzlBwN/WOJoQftCArcdvQwzRGTI30efvSF0f4
GLLMyB1BuXLhHK95ZcdfIdZVOF/sA4+DSSaKWq8lnS34z9yi+mUQdYJpuQv/EBKB
iEhd9T8Wmv31MGottOAaq9MUiqU6EN7jpY632Fa7SflaDpKi5d1NepT2RkarFvoZ
Kb3WZZXONDm+eqw0eE/Z6fviIOLytOWL7rKhVs8h1k1iYnYOUiprVh/6GN1Ee7YH
Mv7SBwix2/4l/a2ik8pdNrLUOhAeLqDwzED1rWwemzgxATTZz4Tt/kR8spCiyXbp
0jZNgORyOgbxXR8k/VkZU6MT3JMvK1Jwng7aqcRE/cfJFBj3U0ZAXD+Tgyg6LuJ1
x+IuyeH4KoOBIzTNFvqt8r+/8Ff0RB+NsOeIOKZ1FbyKue5ZQkPl32bDhTjLulTm
GMbacjJLmgqEfZ5N1Yi2cwFgx3q+3gIQOr+KufcgA3eMJWWpEAdV9942RBovDIfV
LwEsIX2xjrI/C5VnPVIPLwwnknX6yoxuiC64odGFje9170lhzDpkEudVSXXdgONN
BMf0Da+VtE4Wvy/d2H10sPOFxwzsx/fJ/fDsTDHA1kBTvuDKKy1ef0bvllgryvF8
yiisCLjQCjoXCeq7d9yWDh/b7JucWCknl2TT5In2L+oMVa87sSY+HDH3n+9TCzs/
2nOSlxC311O65L8M9XIYofpM8nkzQoHgfTHX6IJN58wD15bosGd5A7GGyiKw9EXU
EZQ2kAopm+tU0i877TU/221HtKc1IioxMjMDfEfVn7lUx0RgnGn5UOIb6Pp4d1yu
d8L7MWX4Orf7eKP0bXCV9aUXMYkg8y3E5h97JGEj/jaxu8ydxt4JgQh5NBw3Od+G
8kHz9n1xlI05maEk+ExdkU7bbGDj0IzGYAFK5tMNR6alyBA/zk3RxAXSqH3kxnTE
g2A5UZ9YjDF5d3e/OAxZ7hRZl31waGRTcR1tMc2oNbKDVZZvAKcF1/zg0TfE7Rvx
d3bquZPO7TrR0SImW50rRVHZxfWTOUlRRpELvkVFq3mJyuABzM1WAbTC7if2b4jh
iy9uuCDXhKWm4Wv7msGr9pt+hAcIROn650KcE8nOP6K7/roDL36Ux3qdgV++rP+n
jgKT+GJFOyYK1xD0gw8Bs8ojoZ28kkqijKgQsLZmAHJSpaZAf+ZDGnvxtQgNchGS
2rloVgYxcQFDERwjvQQeX/SfOeRghujulkVn68O8n75JcnnWLkNrZBo/L7J+0rk1
0vMCSqFClMRdvnXi18P6F0YVYrmn1Oq8r7NQh3ZiUomxYZBvtI788gLiwU9KtVkh
2NxIZxQ1fDpsP3t8VwFW41oOwPwyOSAxKv/AURzDJ8IjKsrdsM5kUQoVehZU1CTj
b5LEmbvtKiSyLbGUhZAoe5Wrz/H/oorTz8mLQL96b2Q4lvJizJAB9Bq/mcqLnLpa
LaNgoMfLsqz18CfdpZAoZ26EZ+7Bcs8TLo/lzbB5gy5p5vLlc3nNlAf6MBx2hFjh
OeNORHIGbBhCDSfw+CWxtbhQQqD7jyM5TKBp5qW5vSP2pdhJw3KJV2Q9fbGsgJqS
2vID9ClC1YlrV68ZOztSyQnuQxKiP0CtXOTf419gMWB+BW2T48r6WQingVdvjuhS
MhecmxmT00dqw9Z0Oa2NYFYaeJt2Ygaj7TAztFn3zAElPi3eMhVx2eu0Z4vfAUb+
VQOTJYA0JlrkpQF/eev4BgQBxXQOVZyG1KOfSv7wVJsFiWu53lYFP4Gprcuagmw7
BbDafy5NslJEJ5Eqs0dNaUS7e0krr7oWLrTapWa9f9S6R6qPYlDWMDISDXN78ZTz
5f+0teoPrdPUOBmm2Q1CIM+lOxZrEBlsbpRhIDdiT9KBQ21JJYEzyAc1ab6yxOjv
N6xgOg8MUwP0PqMlWhsUNLK16wF7sDXJM8q4apof9xHM6oyU9jC0M8zP+0E4D5hW
JVfmX6u082uf4vniNtxgpwN9DbEIod9yw9wTwrvQhUP3b9fflJGH3B/BY05ciloW
nJRZOFsz2p/m3fr+7hRY4YFdOflaP82H9EzVelv790gbEyka4flkn595r1PoIMB2
OZDo/DY3q6KGKtaeuWWvzZtvwjxgASYQttTSBZt0qUtPbSYeN8qCj9jHqJ3fT9Wc
ou/zo0mcqjUU3zjIJ7xEM345ZWDf1yjQZxlqrevLSCxilxITYl+A+7NU0fRAPJZA
C1V421ZNqc7GwwHmVpNdIZpyXDyyMlTWOLLdLny7i8CN4ovEunVwOlvgbYuPBvLX
az73hiBT91+GFQzNMY8VPhDYLqXMARqCdOS1syfu5h9/Q3NyaBmseAT4UTK53Kh9
vBkx5H9CEEjpZDLeXUeZfp66Spj3PQHZRSekvUANUHTVTyuvSisrQ0M5RyIH229y
85aUKLHUf9SvSXePfFtODfTT04vwj3Lk+4Ja1ACPQdDGFNyMaY33OV2vMIhd8JbA
CtTKuR/VSr59Vlq1U+ajQt13+aBDjd7xSYyeYByTfHCYo1vMPbUI31uwU5ih9aag
lCH0QxmfHRQOlv5K81U4p0iojzhcPuMMwJGt1NhzUHsH/VTggDN7mWakpna8/Ki1
37efO4OYzTA7v/SYb1JkgwIdGxewldruCdW20Rcrd+6/IHeqTcpXwNPfTIK6uvOH
Eidzf87RRtxsVKsF7VYw8Aq9HfBUHPPpy2BkhbhkBZ22nvgNchU6lfx+90QK6CqJ
38NjS/ygKWhQ4x9zWLl7T72asXgXY0EjRuDukeE5u4E=
`pragma protect end_protected
