// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
T6O9qy/mPCLrgFOY2bR8GN5l3meAkHAYqHHDTiZ59qr4zwG/WMheV9QbnouNuOVyadDKueslXIoQ
PwUft1pAHqC52M/lX+sZ1KLCKf4AFqAEdC7NTgyuBqVX2gpzIGLjbwwkYlYfjs/bra/y4QbdLDEz
6XKFV/c4XAXPPdsFxaYhPYobxrY+mWZeA6wOilasoEoYUVMCklIEZdMC0ky/8deohfoW2+HX/89d
teMPNZRvuYuby23xBqxohTW1W3b/mjWf9oZrAGUuvt5j6KL6WJ0wCjhNXxU4m+E+CEfHLRkb4hdV
j4JUj/SpvLJ3d8usI34o+gPkR5sdV/mcTpvRwg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7776)
Q1srZ3d5OLr/jiBh/LSU1gOSZ7m8mJZ9/r8uj2HU6NoBmn+53S6Uh+uktU0/WqAZcKeYlvRWeswu
SRa7GrvtoWfWeOCw5AqgMy/5nTqPJ4sJszjBiO51Mo5tOtrzE+ONmspqk6+zJkp7KY2yLj0UQRPZ
OpqeVUGN70rzxbP7Ej7bSbVCfawAzDFF6CaV1kETQbN235ZCrt0GLYaYkPqiVkS+CWNzUAK3r22X
G2go62xDzdsZNS+4kLW6z3VS0zfRrR3PUobYOq6Sd9IsdM3umuYudUt27IP5UR3m+vJHEl3MPlqX
m0FAP/HELp/LtGzA3RskTm1RGfBY7oLexplnZqprgRTu3eDNcXnT727feo0CN+/mFdmy5nU1u6rY
EKNo7Ah4o7aK6YZAtU+CcIC61qghaym0MzX0ZEkInu2x3p7qLHvQEvgIRS23hsKezudf7D75IB2y
/jX0A8oBYXPTpb3iwlKF/tEL5fgD4+ROlSM+/DAFgL+4Y8L2nXsxQ1HKoGFWDBwfzHYVn8kEjpxV
w9N4zjFvZggKHimjTsZw6DMz+FSmRIf9yuPbr3s+wMC9P1SSKmdF0OTrzEmNcys/L6bowzAjEN+3
Sze8mHsgI9b13LOmmmaodA4TqPrlFlbyA6DrhIjxJlcIZEB99fAwdSFz4+4KvGfFzMYe6x0UUQDp
BUDaON/XKsEd0WRXGqSy9sN5WyAXKzQ5OgE3auHNo4ZNh1M5FpXmgSuvtw31pnmuOyhbT625Rhp1
SSov0OljVqQJNtFCcGULGjRHJbyWLNiklnGRX2o51NiJ9fretc4BfOR5rd2PaIw/Cr4U3Au7Bdws
i2XXKfy2ezmY4zBMriruYZmIUx/DhBOXP7D8RN0z8kF/tn73+EIFsrR0XYfDIR4Gc7uGDWYiUKKF
Kr5suEEH/laokHnA16LcbzSed4GDqqoPBJjXpobcEHpMiJYmELRM3QHwjljF9VCe7dUclYIlpQSf
85wm3Sd/6MjXVM2hYJbTgwCJPYFwKomWLGzT1MuYMG3NtROyjbzetudX/N1U/5lWOntQmJ/eixvz
YSRiLqQsWMdJV4A3hYHp+uZtSbdeigxLqh+IiWBb8PC5lGKJ5BZgDvT3LKPD+5ZPd9S/iQ1S1PwP
cn0w8nBQ748vdvPWp/NIJYyEzw2HogUBfRWI8lJ36h3OTRGMyiqgIZiBqH39PvZcEpECE42wXGrX
L6hXAwp/BISRe4n4OC5CoCOwMOZgI1/nu9fcmY7aFBE8GSQr3HFbyK5KdnbU4L3X3/OEBp2VH8Jw
Sn6OnsHOcEQhdx4FlLvbzzGFTyuS/xiY5zuuLDMKkcX7ZefqELnVXBB2FY198h0NJQkRnst+rtd0
I8Tu/vDsSaXnj6l7BEl1VZPr/A5sBDlDWDxS/1JlBMcC/aW46JPgYd59cibM2a7wULKrLbLJSQdO
Mub46uGE74cfB9agrSjW5pDhi5wNhYVScXQsiwsUHAIXydyW1DETa/iUEXZihaSsZFddrqNKikFT
lVZT3eAlR5/7t+JKOLFBLhC0ZmRDszpAa446uLz9vsJPytzBOyhpUHjgI/AzYuvdlXO+EGTOqzgW
jP6fm3/s4f9esDDkAzU9+HYUF88oescb93anRoDSaDEiLCSPjt2sAa3YaKbfRqFYlYo2652Vvc3s
kgpwkkCmoDQTHWEP9SYyRd+qZKFvjvcfvppUVxB0zgGiRG0X/WyQMUcwrh3eI7aRuF1xxfrcWODU
cANy4FF+6beZPbNrmrbWsDuu8z9AE9mf0KXy6UU2bRihH5sbJE6YKZ4DswUXWPM80+ittugN049u
bf+4Z6jJxVMoGX+D1H4rAr4/vv5CJm95L1ZzZav5H/NIS7b6+1kMloOdHGIz+1EXNKVDeVdGwP8q
FOfKpUSbwi1GB2nZbQOCVj4eWVazpW9EDUQeBlY6P7I7ntiR73iBwkhIRh5tT3APqg8WElSS8jPu
gOU90otyuNfY/EfknKrjp0JTxJvunn2GI9aQiv+nrBwOOwewxlIfTlGztUs2g4yPCPdYh8ea1Emh
tG1/ryNELXcNmeZoHHjmp7WAhRXWb/BBbWFbyjxv9OBwR8IWCs3jZOhkn7tr4cRaQ0+ZaEP1dsCh
ffngMOTwB1ko9ypmNhe58aICl4dJlznUfihHgPNcvO4xfc9yUzpylCO0rb4RGodr7TWPe04B2LJ8
qSAWbJVFY0KA0+WMwxh3k6IEwCuJkVBKmvbixuBCZBLzLk7gkbgvGW5uSL0nTN+Owc/CFh6Ym3xZ
jvOKgfM9UChYhedgXh7Y4sEAl6H60fSS7ZUX5hOk6uI4c1GcDq1adaBb41ZQveOGQnf3AnWpi4Sq
pZkZg/VjeymswOf7wbcjRh8/qb7EDHHOWCfIV/20Sgaa10/Cym4PQl1og9jXJtFgbakwRGyHJD0d
nE9tYPI3PTal7/9nPhSXSATIjwDZ4Gh42Ip3+1wbFfCAPm9gJQ1f1A7MxTFg8WyrGN85PwbPZ2n9
4tI8TsQMtB1ufgPDgLdHfIA80EjSpdI4U2tlA3GN3PYf35Mhfgwvtsnh+zQQbdLnCcVZyr9v5wxH
7+FCOq7TF48sgxI49boyHx5yWFgetWaZnnv5pAMcyTaaULd1UdeGHl5BbvUkuqoLN1pTvfHQXgzO
FTDcgOTSF3O1UisReErqtoYKmwU87OvBvwRRfPVFCUPMt2FfuS6cP7I7YdDCQa6xDuwVgRxu5JLH
fpK6vD6LgnAegqoJn5wfeyKZekQWsSRQ+WR3MawLNzyJ9asHTgP1k8MyvWMfPdxWMAdPD8/V9TgU
tE+2BSru2lQnE43Ru9fgE25mZb1Aqmd69WrY57CNAFm80o/d2gIfzwmqljG7iUqA0JMGNr1j3DLO
vULkNcxqXzX0EyFFPpwwFZRccmOaDsQu516l/wYJI6z6YTQn4If3TZu6Yy/LEWo44VNc6hBht+gu
ZIAu4PCJc3HP/ksWrmbD3E8NMFc3qFFQe1FdmBw5vWiMseHYsWwnMcTjmiEmvxzXuxuyvbAg8Dk1
tqxM1WqVD7mJbfWNBywU4DCpKtUmfFYwJbgAGZfqVM9xw5p0lh3iWMUdEHudggpVvzV0cQcplm/H
f41hp3NYrUgntXwKCghdfevhTOd+fREGFGVG5KwRYMJMlfHv3UG5ejE3TJvOakz/PV/PuCQADJm6
Y1u+TDIhhofJqoX9Pej7mqaWsyB0EP+Hti+jhFlenhTybcxCLfm00f3DX3YjmNe1u9vWpJKYTUE+
1+o7izhGeipjozzErqbVYdMzTeOubjWcldzusfeVlpftvkAkNIrHoLmothQ4kjGK8apSev/dlzl0
+xiFg7LbBF4HyoGRXbXXrfBqWh/SkTjTdLTdlb4Ekzr+pvHURoSGr4+RxOfEQo31Qrpvuaqgr6Qs
FFiNBFjqhBgXPjjnSktujs403J6VHOuuE9qfeVt5cKqMlbZuCCqtRSaAKF3DLsDNnj9SOgzSXAHV
PI4bs/grjSvlhE0xGcNEybu5HO83+TR7QGp7gopoWhL+dFjyaE++uuMaaOQ7XlaKcW438FB5bWVh
HRKmvrnhxOEMtZ2z+hiJuH/pCOrqnQRo8BHLrmZIKdRdDUcv7vlum9QKS+5yR79FwPzvjMYVhZMg
wLkmpaDMDm50gWQ8DmyymEYIfs7kAeSqv2EZMzDP9WlOb7/LoCJdqA+hrC8gHNIVB3GM5iXchV2r
Yh6J9RxS4mF407wvzNWnatDfwuO8/vk1p76NeCR/ikzSkMebiTEAzxPymrrURSZr8TebFVcgsvLK
E+Bx3nIFKJIUW2eBl5Dqitsnqy/eoZ7yrn5fwklcts0wkS4TG3IRIZXomjmzpz44cSmc507S8+jX
sxv3SCN3NDWZ3rXXbYunYkRvsR4eNB+lQX2Z25RHhuNKx4Lte3WuTytPNSzfeWkFXmUg05F8iXGW
kVLla8y4qMrcIyFX9XPVlz+qLRexbxb/UoPCjP72VHSNDAbU4LQLmNeN8ZLMx86PxX9f/HmkArGY
5aMavVXs3/KcBub/7ji+ZdcciZxBFQpJmQh/LqtEJ03lB2Ij+SYv5MbCJFaDWLW8jGSVrLt0cx9b
hON2d9LNDGDfOZIR/sznWKy/2WN8UKRKTv8puHkynCrnrbyT/Iexa2CQoiCTyzwsm2jLkiUsPodt
Cpm6GdiZywJj1KeN3zZdRTzmDVyywve/D9GVfhhgfXvJzaUhnKQupbV1XY/YGhMpqcRKYCPjmG6v
WbPpBYrLgZjwmI4xYc19fsBbVX6J0gJPLOhuQCTUZHqrcUiIAdsfX7yhVnpulVY6MbalC9cqXUr5
FMg/m737mZ4GWIvJHXNDkXbGxpwDBJ7fkTkm+PXcsPi1hBgpgpe+JGYGwDqYULaE0b+lsz+TuqHD
d9333pHqJ/ODPfXidyyFOcmt8DwUTAYCikcoRn3LGFpPBX1L/uH9gfINcZxGJOHT3nyLkAkTeh4C
LQz3ezdpwrQzG/2rmiCbMKDl5sKf2sUdnP1/Tr5RXRW0zWOnulyZC+7mDF35csIcAB65Pk1Jjy3m
I0Qx6Pf+FBFvgCkN3H4sXPaemySIOQcBQZ9M31xrFi6f9R3e/lOHKvml5SZpRYhr7+ajY5IFgQAz
jLJG3VTWsRFgU16gZhGxRA6LW1dUetsUUP5Bi3dHpc8VnXEDq7NCidjFQnllmJM8e5gumfZvfkMY
8nptXRLeF7kgFoKL71xRIa6HdaL7aN+BgdArPECRb+Y3/9BokFmvAkYmjmyqUrAt2aTf9UmzJX2A
2muj+Scuu1L4OBzOc6VUDaXVWs6NUXzTGiJr8VDoG9BWaAAuaSTHM84c77VNNNt16et7vcowIaWg
OGUdEQ5UptMETAcwB7gbWUORUH+b7zDal4rleTeOf74gRXeb3iLxWRL+AF7w5pI1KwfcLyGYXTu9
+FVj4lTfm0pHsT320vQiLZzMEASyyOPFSqL3+QFsMkMvgBjHG7UTJJYh+JUtTBA0QaOZUYk83adE
BAAZrnW+6WfsxBycrOiLHr+O9ZE1jRHLJq7toKhsPc8iAauPLUKQul0EgjKg99W5duYqJkheyE+7
J1H1V1U0GGjhC8TW1EEHb4ll5UGKoet/I90izcAxYAOb3ZO7VDRbsCz0DJlbBOpMtaqAXDi4aWjO
03JReKz9HxNz0pDe6/X1zWtn51XUj7OEodKR5mI1Ryu+4DcTk0f2BDiaFKLTQVbfZAEfbnVbdFwq
ZiNrqjPSw3TAGD28pwBTjyUe9lco5IfQx/Br+qRx6WIWdJuHc0mMkymLJsNweEaxZ/8aPkXMivmX
dJS2k/SGIr5vY5hTCebZYBFzL7Od4jTvvYr2yJHOoWDcv2T9luxuXTiPHeBg0NnGWFvY9uML3XEp
hOYB/KO38CwCM0ucWHy5drmUOPMD8onNMkeeJk7CaDK/QKWeI1/6ftaDii+OzqxnUslx0qI9YDPD
WEbageTTeJGc+8jaZELmi9tq7L+nyhnrrlWnq4CGhGmflofm+FP0Q8HEh2zzkYPPadNeH/WHx7Ua
BtlWzqCL0FO9fh4Ah/0TRZmYjhHKpwmiv9p9UbeiwFbkSkV67eWqK6QEIipmZjBShKYOKkg7gIbh
FKNn7jzeVDD0lIPmKKyxOV2jBlGP8AVB69HQmV3XYUYMv4if/5pwYmfGS10d69BI+4v6HgFafUfa
0Ibo+lc/kRQpknpCNR65DAoLSNhiFRM8Y6QxL2pRMwMKEtGI4icVNqkmRqrGKLVxy6lUaEcNYkeM
HP5+ACzKsrvLCOCf3KMkt86IISCACHHA8I2/PNEdY1qewht6R1maJuflTdtpUGWK6GS2e8ouBwl/
dUWv4Cb3Zx3WnnAr3zl9mpUYxUDRV1kmK7RJrS74hMoqoCApNAUWCxPsEpOyCYfTpHX/XXB6lpA4
fzCk28sGr46IIIYIhjfjupaxWVMK3VgqA18+1YBZXdQQKhzqPRo8VwhX/cUk4K+1jh8EyCkVn1w6
qgPGCjATQlg1HeQO7dhh8JWMdfIpdOWUio/kw95EidH76Vij6Iz5/95+bZOIOInuNWMlaD42XDPc
nxscyRbA/VQPg0h0PcDhjnBcsWMWY/ehknpiTpctX2lwCR+LRPF9lTb7C69kF1d1hbmCAsayF5pv
QsLyruxmsQJWD8/DfiW6X1oQkgW1eNxGpVMxfaCetleaqzQ9Yv/km9E30mPw+UWFQ0Bb+7crqfk/
03BIF9cxUgXZkBRTMkmqW8t3RnsltgqU2N3l8g0UO0rye9o9eU1z7K1z+ZPIoHTcAw+W+4bV9riz
2aucYi8J4VlV4shpTV1EpRDemhce9DNWU0dTYhiVyPp6mtiYF+bqavUaNCwvlT2LlbIx6TAUUg2W
fGXrwm649x+e2OMle/SdTth4BduQT7GvqWwR63SXeXPY8sxYn7HNQuZBjP/eEqTrw4GShBa0yztM
C8t9ELhiTrZg1Wpxbwu/zNQtkcXjSdsedqZAGseiTCMYIGpM7663OZSnsLdO6lrL9S0lhdozbAIo
l+ro0bx4LhK9OeJ06wFY6LR1UnVs604TrMeOCkGYItumo/j29zvIqI/iHstxxJxIJ2SKXyBBywWR
Wtd+p3TcaRVmlta3gKxGVea3X12g4ZZK9x8MmunkFox/umFTCatTKJ/wFuguxG6fEnMFltL/gXf1
S9lJ0iXr+W+a3ruCYX7rGS68NpUi3awzYeBEzLzuiqIzzuMBxxPSU7sti6KT9W2ERHF5QU4tzmZu
wzzvKlbfP5GAuERGFcau9yu8nZpByxNVOsZGTg9+SOeQTFHNZJNYaawo6/RWCLQxtld5/N78US+0
WPATgj7acyXA90aLkBKUNFZX3Mjq9C3Y0CtrA3SSXdg7P0CGTB6VD7rgfEbqn3HDLBGn/YHVjL8R
Cjrvl+5zAazXG5AjJ1g3vCxcSvkkA7WSogHBRnUr5o9+NvAPpYOFnLozPUP0Xm+B56oC8BzP4wM0
JOV/DRhk47sdWA96TqN64x4EZAZJIEok1yJ8PMJrUgE6gzSl9E1PActN87Znrq5sqmwxLpukykvZ
ABpCUkewVzlRjsVuYq+QrUoiBa7UCTXy97s2+3xs7C2hmeRxQdFejtubbjOVMH3ipIRwSusMIy05
XKmf/ZCWj4hIp2srv/8Xg6kKqy+vhiZEGiUV44WCdx4DUXbh+q4jk+8LYe0yHgkIMDzbjBVVIg9a
qvw/P4ftkqJDMzdoIbLdwjrJfnVCTxsylIdwj3nKNK4pgrRj1DJsUAH05O18aWLGJtXfs9M+epJ5
aRaO17EnevTtxNlix1S/dc5JBhcgVyHtKvB90AKMVkndTTc0UI7s+5c+w8nMPIBAhtZkwLqGA6wA
nk8c1doFR1W3g3pKwvrKc8I6EW1uB3ix4sZMv4EZUhSFciYq1qc/PvFQNrQM02J3xplATkXC2aoj
cWbxupZsMM1Kb9Oyj+lcQStX+xyrRMwXAlqfCLnKWFrTIZ2fazcK69zHVn8LeKMaPgkYNjUVqlY8
6G6eq5/VN3wdSzwgO8zwGsPyJvlcriE5DcH5ckEkR5JkS4Lg8tPkVWVKBW50ILrtWfAcSge9aYO1
rS/pE3z9Z+EJpYgorggultAK991CGv9orBQCiK8Ck8nRvR+Y7qtRH/HFzyIepcXcoHFL7NwEx5Vs
lTSchz8HciiFqxd17znkzA8KVq37lWhoQXNTKzudMt2sv3bObDcfJqlVLfBFAIjius5Yxpu1vduk
IweuW1BslhawzT3vk0O4g8FmSOhJRis61qfI2olip2eJb+q3KPURyD2XoOfWl0WJfEUexxmYdP6L
/ab5m/PuAJQvLWBb1LDtE1Q0TVAeDXDLsR71+kwUs9f1kKfxI8dJaOvMSMWPA831MN8KYAqUkZTI
HLuT3sshIqRWJQXCHxfqBcfnk3l+Nir9O86abo0vkmj2R1kuQji+OwXiz5dRD8pNwrV5sfs01R0R
o4zhTZi/9fgXPFhDe6ulWFR5ggnuRlQdpG24gpHR7lJv7ycBmojXntrx4nf4DiSyOY4vSaxN+biQ
NX0AId1T5lT+sfi/eA63sRyrLvmX5ksDIgQE+MZ471wlrxzmg4GmoXML2c7Wqco1kKf9YLxEWv/5
qPhkrOhcnbNMaRK3hNKqfHMYelkztYH/naASvg66SplKmzqPUEDBaE8domuAbsvq3EihaFXID8Yt
99hxysjBdttbVMeYzC3Gmo77fgx94XuP2PjAocUZi6ON+Safs2nDnR6DgDgOf7cpXf+JUKw0d6ZE
4gBgmI62nHVzjJJ03UaZAFMaU1FQqARgf0qZfT7egod7epel8j9TCvXrGrf4F4ncKTL2SADfjF8j
1ybEviYOyfKjX4PZeGL9unN65iWMqiQzxPuKLhEcy0M362vhvQZ1UkBBxoZTt1A6xKJw90BUbhvg
2c1AXrQ28IierUFMQ3KeeX7ZhNkdYhgc+i+qB2hN0rBZU10XvC0aSIUvMHlCqeqtf5JomIRRDANQ
mzY1TQolDOrVQC6jHGASaXkScWv0TcaBAojvXfu32Pxv4D7wsGT8zSc160zQFvP2qC2z4WjWNQCI
HbCtLWUe707qaA2BX4PzzHT7Ss5DcgsuHYOKFOk47cS7/3sNrECfKX8vZHsUl4qOB5TqwzxPHl1V
QCtfWSmNWCMowvIcwMDCTvJm8fg8LHzAi0FbgJqbEyiEjwPOmp/f23E64MujPuyRglqPhJQNzKG6
tfgbbPyAr79unyL8VIZ2QDr2M9Y+a+g3qDQYlwRtUAwhdyQWBxPuzJYk/0LWX2Ciq9K6fM9gQ0oL
lLpblDH1W3/uOIatsAg4BL6t6WNHfKr4fE2emNK2ZmOYYxyyzO4T0U+QVj/zm8Uhn8yTmsxME1qB
QNIibQ7TxLmuu/EKj/CuXMXGai6NPSRlwY7V+pePs7vpgfjTBy27ns2ikSota+g6W6JokekvOVgy
df7NrfRmjX66r9E9enJjz7vtTlRw0QUwEjS4MWhRwhOhdgiN4ziwsy8lQHtFB2lmVQrLW2ayV9hS
Fk9W8OQ0JhHGM1Cebix1xOqsIOd8Bb6NXli9Q2OTWTTCRwIrlz28aJmiqpLx8LquHaQS44XrrQ18
XZoWEMcdrDubCSqVoOKLUiRQMfUhJXOOyWP8oCcSoFvP8CUd5kFKWsBqjz6b4J0DAYNK9P6IZbIU
r5Jde63ITjHMMHd8HjJcwbNZyAA/5/jzJm4llfa7KgQhx0VNYOwmzr3EkrBWh3m6bn+ZQAaQosVR
3vTEbyNKyO9EXhUHWiJNhun7co8/lSk/c2HaR3eIIKqCL7+VGZykDoxJXnPwmPh4l7vO/jplzuOV
swCu/5gsCoooXmyC6ZFNIPjhifIpF4O2TSjE5LeT4rVY6POYOZz72lnOsS0DtwDTMqe5C2VTtf1E
zGQh9wIQW2DQVI4cbhpk09bV4Nqsg61YYdCH1+Lgc0enrMIv6Han/qtBmxpXPYfbavvIuqCw3OJZ
BbxaiZygBOnAyucyjdoU7B6skH4M9npKX1X9ktAM7EJUzdrq5eJ++F8d9wepK/wXszTob1z9cpP1
+hIz+HSgJPnFr5s61C7sQUdB/0vi/gxiPDCC/1HaiPYaS0st5q1xhRQWUQ8pWkW45otdgT+7ETrV
xEAZiKiX0K027LO8JJ7DfxR3sJF2zGAXb4uOl/tqQA1IaqjVWwp54mObukylju7xr3AWhpDPHllv
7YmiYoCYDi/XsSlIEIbDurO7S2JwfPxBiKPJysISo9CHiVSsw1EBJoNVWLmVyQ4VpBII7V6j4w0L
yhLqnTNwzcWJxSpIjwCt9O4xHZsUezOi+qq08NHJlmztjTR6eOKvRwEgXYOBFjPcFCVOqi50sPZq
PxkAOTvHfGKlqmtSG0vBbvEparbZHAlXdYaHPkEgoB1NZFps7LYS6kNQAzny/SeZufOQ24ipgM+X
GnbWJYnOt525X7ecv5aJCGprl1jQ488XehWWEx9gym3NkXx2G6Zq1BTtkqufgWoA80npYY0v7DoU
4hwTLah0Bl1YLHQWLvoOHtyD8GW0bv+D9fIk5wAdsrgptp2YFM9/HoEdKfTuYgRh0GRmIlSHoNCu
tNY9vQqSJMDOWtSqlHWASecR0DLrl7Uww0xu/SCeLqSiuV9JDXOvE3eV3bnpP7Bc9QxgmAwOESfI
0Dp/ppD5sxVq4nLFdeeunjmGe4iyaTKtsFLgbNRWrH8O9rqVFFg6/PuV76KeRvnHpN5CwWyZ26xq
5Cd+TQp4x2dnTS+h3GAJz0Yyhdnc+sMDj+Nb7SrsjjyimaY+J9c9gRle9BSRhusUHdXWDanDPQE9
fuQvBdppzFAqFNVk2dotTj5lU8esvFJ1
`pragma protect end_protected
