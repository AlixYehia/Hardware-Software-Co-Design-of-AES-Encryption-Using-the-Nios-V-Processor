// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
bF/cvO35RHcycfec3Y4pA+GD8iGbvYgrZc7vA+1Mv4PR7Vt2zheD9/lCoo2FSHQPSx41wofi3uDm
DT7IxMNb/y6/lDwdVUE9BZ/ka6rtr/BPfwsi6KkoQ6HKfjFSPcVDtqg4nHLjbConcQaKlnW4WzL3
VEFC54LzNEr7crEAKRNZpn5Z89lf/+BVD0WcUAoKX9z0OWyDxMSQuqda9gL+YcIKe6yEg+17Offc
3kMtv2Notb/HuhYG5GWGerFSvCVNtwMfoUNUx0R0Ir8CLjfrPZ8SqUs0mR8nm5oaRUoWkcF7TNkv
NNnW0tef/96yQVeTyss2pxlsR2JgBAM64N3BGg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5600)
OhAjixh8gBcdMDzqsQPZccs1T5Gvmpu6BkrY7q4CJTOfglQM7FAu56R8weC9xAyosQtCp6hHaaqN
xlRZY09202Kr3laQb+WNHLZMkzp5wrIWLBoidpkhterOBAuFnlV1afMXAvK1J3WsZUIKNEFRyUUa
iK4v6k/xAWJTabXKA6zmlte4s+VR4AP0F5GK3hbVelE1pUBjaMneji9HvmPs3FCx4AazRHpdI92A
K3S6cTCuAKh7QbhhibwutisfXF7jIyIqGYjy/InLuA+ijyWraQGyZnnGTb5Q7IIGMnPm0HSHjb8O
SXGR3JklA4IFnwx6SZzDF+YwQnoZAN5+eQRlYdOuHqG0Ju4qwpy1OaYyD3+hXA4FvDjkcu4jQNZ/
Dt4pKpBQRLYNnTSOqvyY8QLpacJx083ytL7tkE9GYUEoMB63VBf+cfC8DnlxBuH0fHjalJsi4Zz4
oTePR3UrkgDMvw5K3b9ukshyr2sLeF4sp4VEDMSmQ1CT8lhyBAp7woBFQ1cvAQYKAN+2wNY8dAbT
DSWvS3nH1L5+N/Zf1dOsKFiITLDtg1bbwsAxLjRNOeL9N7oXhGBb3UuxozzjLDpG7aAtIm47Q+KM
dt+bZ/LEyCr3XKMdKK3+xOATzD1YiBGQu356ggzyTAIldM0ldR/+XPOTA0VbhKr0Jgibqntj9+5B
hNuSWpdHWH69G0YlebcibteJj5bGO8PhdEaRTiETTjftcbJ0HOcI6s5doBKQF93UhwHMUXliupzO
VqgnVCz1PtWztkpdx2DoJf1KD9nlS2c2eY3o1tTBs7So6IiHUKelHxzcMUlqhwyhi0mTR9Kg/nt8
9v4TWDro0nngKS8j9WdgXqhH10gLdqQ85sxjVDIQGotDCBc6QQ4+T4wRvFhmJGNcAl5ZB6WDlJfE
X60tJ78jqvAVSb5dZ6WL61rTVNzmX29AJubpzLxMhzF1CWcIS8ayYDKPXaSe9DkLLLtRCpqR/rRL
DgJ9h/PWfdGrwXr4vCdl49nGL69EJE6w6cvkdGr6j2lMdWYkUgZWjHk7kXC6rfiVV+WnKZCxOk0P
yKsMSTuw0/kxqXXiHt0VdS7h+jF1+B7sZczLt5Gx04s5gJpHZC9GlgLgpkflSOPLC67RjKY+t4k3
9POqm2IMAIZL+pewNOw16xgwaP6VQ6RDdtvv+ZONgwTc5n3UAINrC5kTJWPEQP4zNJQmHMvnICQA
H4PSaLo3UAKSTaNp+DtwiNzILy4/9DD3c8b4vMCZxd8d5uYlnvJ3Au8hTNXoWS+rJUKKRJU7ECQm
7wgp23idhoJnSNtXQx9xJcVpha4p/nKbdaa8w5GEVS+Bycm3/GJXPjz0RJ4V7NLx0MFFZxgtqAKJ
oa4TDlRd/GKzl8ySsyJzO5mYTjhyJ+8dY+HCUEtz0e115PCjnl1Lo5JsKTsytXyKHovjaWe34ePz
1DoUhqxkYfiWxxsSboFxgp805ffJ3/TuICqNemwrhIWq3OSmR4hkyD0R9tFGoIZDj0/pSrEFgM0D
Op2A/Nujh3xXtPC1Q3lnpq+4O3iuzVaH2Sv6cZP7QoF7kdw0K0wpBXKncWvir4B9U45u1m9xEtZ/
EsQ49Cnj950VuNhppMruapRgryZacR9Cya3PxL53KOSYQbSiKzZFQqnvV6OtoQXmt0f6jqnEECy4
gfD1boNexdCkV9A0XqHuKbh9wg8JdMDjQT6bhWlxj7fhB3PVpRUOJtNcOzarncVfcJTdVVQcplC5
sZbQWvwe18afGaSwgSW8TW/k5AwlGq79qf3DooBzTEaeBAJfjW3P/Qc3Wp5nN09pjdm76JGeWCvA
fMMAA6IUQLmAoTyyAHutUVqaTO5V7qnNcA7D6iO3tje38DEx2xHQAG1Ct5Yx7w2Qn0Pa8paXIQrh
JiFghsSmi1FYyLBEpLTbeC6CUQCT9jlVxFSFTySiSF13xpLI/+hwLyAk1jx5USkRkmMftNFvH4Ax
wv5LRL9KPBfn4oMeh/HL1kVno9hPvksKuhS2ascUxkCXIIm8VYu4IhicKPqOu3Zt4ecmslhoqwF8
d+y+lyNT6f0T8xCZkQ/aKNTpwChq964iF6NHqaieF/omtkL84CPq6IElz8DCQzEqwGMlTAXlmfNM
Ec6rAQ4vmJHGtYI49raTcbzu7OSwc3WdmhrTFdBdD++t56YGPjvr1L0RayGMfZQ+iacWRXMevwk8
jsUq101q2syhRBHhj1BtCXnLd76uD8FgCjiyaQZbWV/lzHGd4NGq8kQu1gxyYmtHODCpznn7VpWp
KJm7PWZ1Y6MlK6krTWzpEW/Fk5RyHFrog+/Lj8oXCkyp16M3BBsZ5i8XRZzxw7608TWvidpjmaoP
5RJ/4dpf2+lQO6EO9aIzOeox0bARwNnZ/ztoX63buBXTW/vcDiG30fvselNKTq5t4TYnet72g8YQ
0RvZQN8sMPmfvt4A2A92Uxy0bO8wkXuf+YEwYWv9/1TMsjvVRjt6hizQlR8Zzq2tryeMUoNPyhHI
lZACJVKKpkFrVO9xe/AkrifQU6kBYzrZcW4FHlLGXt1Db7FlBbRJwNzaakVLVu55hxNS1QxbRTbH
E6jZgi5qKiOvhDIj/uMFD4/dgK8d1nDQz8mK8E4YtHTYPhSTHgKhezmpQ7nV+nCFuuUYP5Q4Xx7i
SntDIaTDVmP9Xue2cxnj6ibJu/55/PTOyJMH+WuP1c74KvgkYGUh6X8aqjG97yERQiZOnknGXhVD
bSQb8RtT83h+6UBvxuB/wyEc0FbnsA9rV0DXy8KnHLpVH1fYDz1507SyeqmVLDAPxPbQzudlPXoE
qjAMY+bsD/2YHXU9DR0b7Sele9BTdzj3f4NLNrFR7fw42nl80TccGg9J0wP96GbeOsxpGGo1qh2p
G4m3SkxN7nWUtPGBB6jYt3VcJj1ky1eAbKAd98/AN15uzoTo7meSahwSsbFbfgKScr+6gBe5pBrE
QHnZGeCV05KxVZAG18GcvNVT/76vJlmlyrywB6mVOdBf7knqVYHPCrnlxyJhOoCLsABvTgVASUii
FAeLaJJMf/hS7T58zCA9cEvdrdoCttzgmAPpdmXhlBjPzGsI0Eu5Cf86j5bte4SqXp/bMolJqEB9
xYYSFG5FnxyuhK1oUee6SHrEnbBEsx+bF/8aSaVjPcbj7veDnSE+bvLZqbaE/rgoNuKI7JNDonFT
w+Y9xrrwwTOsXH7EVlcUx88mFLY4SwskoC66HwWrkEtwRnL9NjL37q7+mLOZKqBO3dxRwlSubKaT
UaPRAMg+c4ePmTBtHsy1TDrvVvq/rgEtwvnwZiPSk7KXpNZubIv0JAgVYYahv98sl7XNpT1+x6ty
jvcEjpBuiY9JsU+hBE4Whj76DcmCbVinimU9EpD+aPLLcx5SecTOr/pRROiunkakSMLuGXqBSl8v
QztLU74weEebiPfpDazu+HX+WHQDzllaYGWQgWJ/+Q69vPm2vnNmkoBU1rIMuDiJ9wYNl0SDOZv5
dOWIcCqBD2STdqjMqu8/CYNWmziW3syoWRhZLH7ybLCJ9q7pviOyAVSLi/OoZZprWxNFjCWqSFK7
zc0AXtpfPPxw+FNBWb4m+xK833vJ+HDIV7rFDoJDanGkGtNMaRaxHheobCoNgBEbzOTxZGFMo8/l
TSoBtBVfharoSrWX2i+9tOKMremTWMFVZHTW4JKHMwBLC4zs7kfCZLTdNsAPZfGMC5pLsQ3GEjAK
wnpF5Ihwnw2EWfS+ZmHTrBmoOGfc0LyM4TZnMihMQw/DQJOnzRlTFBVuq4kRg/j9LB9cCxLarx1c
aQiNFmNwVctPEWIwhMQczkbpdI/AVhXJW+dlJM56HS+a0yvX0LZZGjSTGb+7vNImuBtgkEO1j15F
naE/FfpEDDOud3rJDzZVz8+GjERLEyKB2NeN2wH0MTzp3HrJVVwFU0b0ocHNTV6+utx5E/ZeGQLb
ItGfQyltaJf2iPRd8gVyYDqyg1x/54w9B3teBcDSt94B3hkASu+k40RbgJD9P+dW2wMxrVhCdr94
ImyXnmW64qxDbZ/8BhKKShEaCAx28ns2yM9C9un5J8Y3JVQHtpmyBY8xbUJAPBQFrRH/pcsUkdid
XkjkjHf+vPMRhVpRi77Elx51e31QE5t+7FIuBNkYMCXNz3nP/CE7eDtePWbRKy1IK5aHlQMS2dj1
EHKow8xV7HvBrTtUQ3FoT7m7Ld2uuWy5EKNh3M4FThuEDcuOR38/12Yt/7xjqygZvetn7pnOgQY7
53acLjV15WrAp10qmq1xciU+ZdvPPaxnSXVlcHy+tTvvTYYh7YbOHXeHFRUMBJd1kX4mx7Ng+UFq
p5gYavP4pLPV2Q/BT7F2whqwNhC/cG/NilgV8FPvNh5nsQdHEn9eKdPCfORfui0b3LR/UC7S0Mt2
ECl6c7fzEClPI3KNd5s4bZSkQ9w2ZJ+pQJBcEuysIxevbVV65+qFfstQH4hovc6QjgsvSklrvk9R
Gw/q6SmTlcqJoX3cSeBY5adlNPREQAgOnIlXqfszbpEn0bbbJdL9jZGt6jKaRsdJNV5yUVs+6OHm
er1eydhaTEbME3faOQfdvXwssanIo+H80qKDqjXAl2QckQugG+4Opnu4c5vjqe04rFkrqMBFt0kN
RmLCtPjjp/M73jHipZh5dNT704tPhD5IS28NWLrfugxZb9Qcs72MyGiN1DVO6OmHGGlg2w9XVVDC
mB7UYmDHPVzCPKLWaIBWOL+vB6EbvtpmCSJ+GofV0lxbGOWNeEx7BA5X58h+puNre9M+Cn7kkzeN
+ZKOJHH+X9Hgka20AS5TXrrUxCVL22lxi2R1TBEPZeas5Yjt7Nm8HhJjEoX8LD2XPChJ+eJ1kd9K
wPWUtPB7kz+2tODwxim2AD62dAgM1JLn7MaIanMbf1fXyzPgMb72+QtFHys3BtmzPJLamyihirvU
T4H7pgizxlIQoAMDgR2w7u17Xu3QVlBJu88mDlSEVUSAqskUSiXxVfUYm98Nqf0tejOWecwnJWcX
0XyVr+h6hN7YfACXBc8pvdG/qefxuw5gec/w21fD5pONoTt1X9bbHEmyPOMAGk7fmAlAueRUPpre
opk7bZbqx8a+NyyFyGNpkkNG1kza7Fp/ZSd/w+O7ejn5pda32vLrgut3h27j/0q8mM+8jplCBMOc
r+t9sKJGRSsByMbicO/r8CGhoPD+Y+UShC9bP/O3EyED+QBC7Qw06j3UlnjO78Jm6uxrXS7qYS70
aucH3cDGXG8OCxcQ4if9RMrOsKo0Ga5QsvnWWSeRgSosMP4ronpo/vwqNFx/qodXbuHFRlc7TzeF
HjmNqKIA+rAUA/KBUi65nO7LhMgrkPHqQEE+H4hCJ9RdwQQ0eUAs9IJa994sZFi2qEESMxX+PbHO
otWtwgkcC17rnlHX7gCrPhBZq9iHKjUkU2Y+ds1js9PTfRMGcXWcdRnk8/g1qXca8CKyVvL2ee86
cV76QxhJj3VXynBwYxnj1jjlaI6oBlnGsS+vh4+F8Sl/tahJb/ZDbmmfyR6WHbn1sThxjybitsv2
MfKE9d0K3O0zcn0nj4L0BR2DV/nEa3pL1zYW4AMHwMZGp0WPs8ChNnzsEfNrALBv06PNUh3X40ww
Qe1DDrb1wm9bFG6cPfBrqHtHavIi2Sna6KEm5XKGnAL4AQcWoA3/eX1LgoqqXjyyXAWgYIdGGxsE
KUZnZjKvP4ib+EilcGj29663ntInHDFStFNqM4fZSWcMsi3wjzA00R1Ff144BDgZRDiYp+c++u+i
x5lw4Exaz2UxhmId1PLX6oXMt5QAe81GCB1LBfeGlNcmwVwEbZolihY3Qzo8NAUy1F8HG3LgGoNl
oYkGoYOxhAVbp1R87u9m2X4RwHwy2XxuzflXhNo40iYE9UrxzZBhugzXxFcONuROxI7SGzgauvEJ
p1pAcmXdFRjlEEMa0QMkFtoSn7l57y3XuTSEUgTXPmK9GaEA6i3DuNAp5Y3cVVlxsIRsXMGlu/bs
zeR2ngPTiIBJVWGD3w0oUGlNm0NIQjpwCzvogZYWjB1mjhKeVou9ACqc/kDVEFGD9Ra1lEx9V9ve
7Oltr33edhz2uTLZJmYFXfoj8mBfPyR6OaYgZ4Kk/PEqjJkxHRe+5z4Az+QVspdr/nPM8EOZKYwK
EXt7p8WFM4IdafHE3Kzna/8nAl91LDVUtWUW1IIn6mcW0ZB5Nt2JcSie7mM+CQODJTpx3lbLZRuZ
mblIbwxhlbITv6MoGyUbAQ5Cfvlh/gLpWGFW+xMc3LdgSFpUzLG3dpYjNmgAS5do4abzLmFAKe7a
9oH2mgKUjUarGu5wcafLoff9P+ytU8Iguv6H3b4PlWgm8dr6svzTkVjnZytBPiG0JQKSuNYUzM/U
blW3PSsgZEbK4dxhEwjVjkK2G1Z/nbs1zVWR1yCq2/RtqJ1bcIYn6RM7BW6w1mGCN5nSCDEG2ivr
yP6gJlQt4FsNtrnoijBnv+oqqX0ZkxMPoOGnMgU93mueC8S7u4HzhQEloapzONmCUMu9znCk5hEE
7N+V6xg+oKD4q0MM2f1bQTVaQytK8AH4QTyGqpEEKg6gkakyipHcW0aetoGJrxL1+0TF8VtkU2f1
Th3GT2yp7diXY3mi5TWZgSo5uXR2yipPEFVXi8duKUHwjf0d7tDgIl44EWTp7mIr22SkJ89owrxI
+Nu6BoqGm7X3qGsAQ6Z6WNHqBmbyPEDov5lBosXrNUUHFOMvivd940YSzUyCpTh+dDeBsRDNagke
+0xggT5UUn5mMRdIfhHo/UmLcO71IvCy/Pkn89zu1Ucjv9iQFSbvFQC+a5DvWom3w7g3k2wwzzBY
mBdva52BsyDcCfodrYgYiQvmy5ipfCh3VTN6IMu+U91Oh3Uf4GJR3tcEpPaSWiZOaA64bLEBFI14
5wpwza7fXcWIBWWCc/EWIG4Rn26gbfQXyGfFhKJgck+LJ73zdkyuCCqWRx5chBhkhBsTKnICnaIB
R5S1JM0kuWtXms3PdAA9cSjMsQHY8NyIo4G5XIekRd4UbrCWZ4oY9uio2rmzjHfvjIlbKPpOEPXh
u3Om5TIQRnOFkYEQ/NkGMtA3NZT/rKjI5zXNAfPKcwzOSoKk89QEqr9JbHhD81TZlFhpKrSpLzwN
cjJevt6DOesAoHjivOOh1RAULp9UzElY+piBtPbq0uyuP7+QaT6ZZEMR4zBO4l7MjGTeUcMBimFL
GiZVo/WVfOujFggR4penV6DxPQt1Q8iKNTxSvdK3ZnXqozPq6hb5RbadlxDahslnZhskGYIvidKh
4U6pvQGFJaFMyvaFJQcbJApOg02TKSakhCxSE4zNZsI9GNbDsUKrAWMCN8IolRNAT9kQIy7l8ynC
IGO1mY/rPwWfA4NmkV+YplZ/qUJCTl4DGfxNV4C6MQ0lWyAQuF0cStl/HDWH8miOVCJhW9RPp/6w
VRFEwaw95UEAxnikkhM=
`pragma protect end_protected
