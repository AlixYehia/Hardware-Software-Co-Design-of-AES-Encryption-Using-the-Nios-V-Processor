// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
YyG02S720ZvKOUxSRReXDaqUNRvpugLkbo1Gs6vOf8SLCTXzzAM6HBonIxuv70ZUOWfx/AKYXcJK
Fbwx4iwgejHE9WSBX2YHiaILWq1rG5VIBoh0NN+HVtwCVQwuKNORBoAwapeEDXxs1+MJMzR3hXpD
TvlQTgwgt9dn3to1ufI5LnnV52BiRMAdLgrGvRdHcUXqDH2REgCHooutxgu74w2dDf3BT5liiwtP
5zvv3s+kc8VTCnvagNn3fE21OFjYRfNiydDShgKiPzJadjuvBIVVm2s5Xnng4uhGBr6ZtO1FYSRX
RnxJPER65IAs2X3HsB2DdV0qK66c26aviK5gqA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2160)
qfgMTQzT6RvQE394W8jQ/Yp91RPRBVhrrHFe1S173HMgKXDw42xFf8VZyW7QBh9fw93eAW4WOM3l
eUCtEloNVVmhgZq7rgjwtaZoRW44FjmlXr8tYE6O/udh2mGG4EkXDIF5xVa4cVByOn1eW8+G+KxF
BdrKIArmwt7PcJVaOwAf8rVzrfqYJJTyfKypCuzEKkZIleHVjhSewLkBk7I6hHP0LNAooUXDuPgL
s2GKZ69nZOfdR0tzbqU2UFTtUCV2ncia7WNWzD59bGOsqXkutOO9/y8kyF4QNZOhaxTuMakTsxpQ
pJ84E8QzSSlIrSdxj+U+0UnAOD6NcYoRr93JoikiJDHT47eVbn+P7O4tpS184BzoQflSJ9p6kV+g
pyp1EXfWTpOImSfNF2wSWxmotx3/uW3ymOxKBjn1ntvqsp55PYydmLy1wcvzFVB5EX2pyj2N6U+0
xZY4p0ciAH3sBigw6rd9awO/PNlVrV9z7xnC4TrnT4TUyYmqshuvUKQnDFzOSeuMFCWfIKp2caYW
y4x3yE3yEJ1a+wkaE7a3yokzL1Jl1B1NwpUVvwWQEMBdub9AgFODLbEaANG7VT2Ewd+dRCPd4zof
NdOfu9fzEZAb99qyXeGQAjJbzMN6AaXwRWcrV/z54O3UEdp8bkiB3kEp0PEsby2+6eDVOhPZ8Ac+
S0QT/E0894QBQTQ16lF9NGbnIG1GGEcTxMsPiiOSJgZwQhx0YBv+zuVgYM5ZBfcCdX1dECt5iFOq
tp1Lrq8vTfCv+52lx+3pF4l23/QxE25JGsRM4h601E4TXNVqy+TQ2XIcLE4u9Pb5lvGv9iS9zy5X
WNg3CkENz/+Y6Bgn4LPmCeK5Vib5u5TzzXWsxqbVYzyPU+oORPWY9K8iGdtkxcQ9YyijdnKQAI9n
P6tmjm8BCCHmSbsaFInCdxlhdhhlP7oBfj1JvcXyTQYuVFw5kzraIR3FpGkoLhZQKfKyHQMePG3h
AZxTX8pzcjV/c1LrDTTok4mDTWLXia3V2EPzAuHat5jGtX/w5Pi3D3aVWUqgG0h47ftrewnP6zD3
K+eikKBakE/9U2w1Ji75ya+Q6J70zYA184tz/qJtfsZSEsVz9P89qSZJp49xPBdRSUh3lvPJV42l
He5cbOToXk+8iqZThtxlGp/U99YUpYXk8gAbzPqDdz7XBe3e23/+49Ec5kbbTEU5aqvEALXqhF00
eUm6RElt0nAbfQI70sxhbcxBAMQ0po6cyDN3m0kR84RPjAvcJdqr+IIoWHerVug/AsKrBZKSG5qn
pCneoEOoWV6Qw/zGVFXGLaBJa3LX+n3q8CuyifP8J2qoM0VgwOHPNf8mGQ9MSZCDIrv9EFPdk0WT
GhGMg5bWMOqa11/iZr273OOnTzMMHCzGZ7V3e/m9jzlDMl0YaPO4UuSikQ6V0H1Cf5bk+LDyX3MU
Yfaz31p1WNw/qhBeEK/CuRSmJz0Tk0iAB0Q+pLMoPtS7nINdRN/WO807araD8wz1/8ydLnXvRZeL
w9+9roFAHBwGMphNRqfMjjXk3A6mbFQ6DBZwlmBmIFVVMz4Qqg5MAHrURpEBsSlasvxAS8L/HW7H
Vt7QFRZrtziQTLV1ZdLv2PCByWa1QHLlrew9b/9v8847xsAOtEGkyMx2z7Amlc3BX1Lr9YsgJK2J
TuRdpm7BgMVqexmFm1FZnLPqeU1cnKi1OFHiHIoRz/747MRDncPzN9/PcI9GP5WNwi57QCfjD9sC
VKjDQwEkkTeZJROhFvJf1deTvvvOwM26qm/kg3ua4dxstDMPXHiEYAkRk13jijZVjOUH5Tve3JAF
UiJaKrojaK3/W9DMxxv+ISuIOWFliKNcCOKNi47ZEjyLfwk8+RTdSNqbRva6MyKtIFu2TQn2htzJ
TMvTt88aEnemAOF+ebIGYJr1wuP5GQnl5QIfTK11ahnvRytrpuhlTBZa9XAwRwUnBLNRQ6UQIxHR
TkmHZ4UmTDLs9ugLjcSaiPjIGVf4PqdWj1KDJpyUIbXuBAMKPS31SK+OGSFiZMv4BDGJaUf1zbDv
ThlIJfs7HFBlYCLmT4cmBInP/WNURz4/hfwOhDPYyeyyX70k6JGh8BrSiTC3Xw1tQVAyQWrjlGsd
ZpTGYQJUWXs6uNjzog1r9+iSmRlYpvHgZF5OzMqMGRPTsdpL0TVT9hKrpZotLCe7uBwDeBXUJPiS
dgNMHNzICieaq+czW8c+7PwjoHMQkZUYKFKE8FRoPuJldcKUWhOfC8qCAnAVX+EhaB7cUZJO+ktT
Icq61R9wwC0CtwXV4qO9QiyeMq5BXfseq0X9yrs1pdzcT+49nRh8bFocEAv/XHXU5YC0A+SdUgB1
U5BcIhSMaXVofLGFbvBf5T2tTxVKtK0ij9X2eWfd4Z8Lq+cCl5yW9BGwiFvRs3wRJcfrNqnAfk61
iPNqOnhVIIycqxoRpjfJ9/jcO55VVsyPTVFqcMbX5PwTOhT2ycU7Q+bCecFUfjmiJ8Fmx3NyQmJu
lL11QvDrMtJkZbiwfuz0GdRpeCglp4+SqbS9Gd42iaQ85GkoqrJuoPk1R0D3tNpoTp36A7fEBxyH
Qte1wULRjHB26gYhbs8HeW+yguakxAgHifWj0xJuj5mY3EFwQZ9b9CdxcXo/KOOAm+8yd+D0Scrr
uq+CmRu0U+6ga3TIm52mnVLbeXG0KTeRiZxN+Z/MUfRs1UqHUVSw3W5+HtTWTy4LU6/4JVWc0C9x
JNibsQOi/A5AFGEFnofwSVH9hGZdhfgQOFLqbwVwQkrTu3FchNIIoise+9vAEZAk/qKoqUj+HSTj
Lah31YQ8XYviM3hcuUHPeMi0pHjkkBgMUjs0j8OZ8j/vJvBCj7R5qH+bd7VjC+4G+yOd
`pragma protect end_protected
