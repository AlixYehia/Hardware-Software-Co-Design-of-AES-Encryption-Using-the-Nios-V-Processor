// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
IBx1kZKp0gv0hm9UDLP3Yhyd8y1JkR6Y3eSzTHiAUKPlNhMnb+6V/WTA+HVHE6v8B8fM5uh9bq5c
nAyNIvMSkQXVpL7/jkbbT+iKnUN9vxA7TVgO3H66fhPOFTVbglL2weKyQKr/KTif5d85SuiYWP0A
aU5demIuDaBCyIKWxrxqYjWIYL0Yn8o2WtOjjDKFVvSe12/p67LDuzyML4pD43TgCBoegBo+kJvU
fvDSymqjjhV3Z7Q34X1VtYNzFKEzes3KbmHhxBXtAwBGICrefUk1ShP/4tV25hVbjafvFv0yCdQW
og1ZBKEKm2Qx27BK0iMMGyAuu5PMOWh/tSuRTQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11904)
p4JBEFemNEBK89tPmNAJJX5TeNQd/cJ2TzDaPttkqcSJtN3THZYBq+vs4Etv53LzlC09h6ZNVlJr
ZH9yB0zkg6QypmqkkkPfgWXv9YuQqGn8NoYveB8Rh/WXHGUitrsRSXnRcOyIfBDd6FWT7izBYy+W
RIqtvYwjJq2K5Jm1/NIRvPKbx1B5kFBiQnD21kiy1IoApKZkLhEw+59LzNjr3E/UCb15hY2iEeXp
JqTprtmWvzMCK7cIaoNcveOu47PAg199iFHT931niwbUm67qQYwZf1iXayDwRIczVBoHyW7+lPD/
TOnvzVrEGDOzh2+Grlttc0L7hI5AB9r0qrM4k951/W5TSPq9ZGh6EW5+jtxyqU7aAi6ipSQkTN7l
+VYXfowU/oe2LkUGeslC1bHG7n07dfmEm7Gfl+XjyBEemDQUyfErsGuJMGOMk0sSQb1/wwn/tKYw
awJf0efvwVlHSO9SXPLpHztj0bgRNeQ8hP/1p0YDvu499n/4YWII84C4G0szaIiZhHRkWMbojeFM
g7JFsYaPj+rDu9QhQR2D5GL+MNSKDCiyZiUkuz4ZwejMGJpoIn2RzdeQruWiHFdsFx6N27kwPbxf
+9xksHuEipCMaayOSAZypluimLUNX0GB2n3iNRAN2+AB4AZt3V8NbLZSNm8zrJIJPkCZIbDARZR9
RrllejTDzvXDgF+4WjCVx1ioCi4e0o7ndavun0RV33HVLIW3StortHaFH1j8Cul7PBezAGPLLlLg
Kojes4FMHhvkr1ZMO2JCtisszOajlWRBStMhDWU+ga+Am95Zg26Mm9VZuPa9K9jaeacLATEL7sUe
0nvEsOtyf36eRY0Z5McxiweZawK9itVs02tuOJwQAE5CMldSqhOJhVNlZAFR5djqvbmil38pVk/y
8gkf5Pj6XpaFPuOTQEXMMLfpbcDstv7DJwIW2Y369A4v9dQrCIbbThLICPXw2jDprl1NY1aDE8d/
SHaKZ8Lw8YBx3zyAMKE19feRpK02kiG740JPfGmH4OiGyOeUjmr1MQ/cAk4Ae99moiczBctqKoE1
objl7hmkgf+Zv19dDgiemCN1CSMgAu/9G7sfSX2f72IZ3kUwxFGsdOMp+nPwyyg5G5hv8I2uru0x
36NrrQaDkB0ulFt/ffCLE9CSg8vcdlJR/QneceLqKQBJWzoN8Gsr0+CA/6mVQ7dsPb+8c2fBQpQQ
FnfhipW7BUaoOTGZuVHB8t0EdJ2ObhCliMg024tqXEkWGiahPgx+RdDiTpBhWHlMuZ91CUD1SbvD
T352lKCVc0Zu6fyQmvu4trj4kW2F5PRxSCh8XU+SQcTwgLe1Kg6SiU59jz+iZlwRQ90IfvNz+vvH
aT99j+NTekEsLo+VWOFDtc5MdpyJxK2aN6Y//yDKn6GlzTv4xB+civ6G4dbHpJTzfWCYpGq7oZml
k+UD/IP9Pb8zdydAo97nGCk2xkaxXIHe/kmyfzLkeY7n96pFJyS9gPrEwsiCUR/Ru8a6ITbxh3ol
dbxyqoeGI6lMEtuFGH1Ki3KZxxWg8GjvCO+AQk8jYoTybeLnkAiT5Q0Mx8b5+2dVP8fDvMDZbTKc
+Pl0V3QuD5VhEw+uWI9uQolKP9Msc0cfGAYnGmAA8VWycHbjHNYAm/9tYmHUwM8lQ6/7TmQzOJV6
4kaHdtLazusbe0e6guVPsJW/xSygJoQkhiMWxjmJkkDne75UPvF4tWXYDEBAami7+pepDtx9KZxW
WsN/Gdwp0bCUKX9q7C6lUTUew2jRWalq9qFJC4exmLMTwajAuowwcxeg+NK1e3ZYcXT9NqmxKFbn
HhGve+cNBhrb0nh8KM8K1wuJgmLy23Xb9FepSGvqtnkukwbQaq4IhylIwS2A/6VHm/t9190y9zzU
wNBvmpm5lMCf8BKoUfYMcqlGJ+40e86rBJAidSuRkMF+xIrtCl5nzjT6dmODj7rCNB2uQQhrqpvq
pug4HrxfMjf5zrwbO6WxUZt34xsMVanekV3kM35G9KMb0hlH3GTX9JjbBya/wGghdY70OxmZiKHJ
CinpwT3wo8Q16plk2Xm5nhNMBOi3e/8I4AZc8CNd88Rljic7YhWD5ak9kKORKhBkldbPxP1Zvcrf
wf5+ppuY8UvUATkFYrPbJJku+mDoLbfO1pbkpUN/LdfLey+DkJtXd+RgS6jn/rQcE6iy5R/n6jQX
QXnNZRtwl+agfRbXNTeFVFZk0x6Pr8KqRTOILkoo133SiNnJ/9hfuLduxcAXcwWfKusZ9igKxk7k
UYqcIF4f5Qn10uiNAcv1pKhgvqUWOY2052OWGiIDKPSl5LWNRkhwQ/XP+Ttk3/5NFVlnsWgHQEnO
30HnXCoqfcHlsJ1zW4MoltAjK6QmmvgDVN1hAYYX3DsCXVQuEWPhhkt3yJIWjx7al1Jc6wvbQTy9
prEzUZvRrmNoPHvX9SBQSG4dY3BQfct12kSP19Z2OJygBRzZzlSGHHGD8lNZa25fupal96LxjkTd
NJ3FIyU8VR1Dd75A4UP9NSIR6ePToeELLXf18rSbQVxkoO8R7mhjIz0jWXYlZV5KhV42TLDlVH0l
q5fHcfUY0x+zFnZdR5S3eMvvw/dZ2h6YmdNG8EedQGnVc0bJPxpVYxK1S8mX2da5nQ0+tuGDsNpJ
YSfwDCOq7kKJMzVYS9un7RhVhwPzvmgEY4OVpLeIiSW0IRAQ0qFmJFvz/+Qam0otyC/tVavgq9fy
sF/qQqYylNcnGHyIZcxryOx+K+VlJmCw4k+tQ0JOEElGyqXxKGvLOoK4P6dVU4BArKW2Tvm7n8Ph
XdhUPJfp1ruRJHwM8uQ2RI4v5+NO1E7EsRLIub6tddlcZ+UcL5L7a+RBqrk6Mc/S0vLADWNOCFrg
5fzsA/TEX1XvKAGtqnfjCioBbxBECBQnQTm4FwmsjrexaAYjtDd8wHjzXlsu1szA8ynZcg418B4N
nUibB+DdBDXWv3OYz16wiKR1IsKAcQmYodDi2tiqYsL15mLwDNQ3tj6imOGMmc/lGl89uDnRaIuP
w/sXkmVqSqOJ9mSqBJKho3gGjt9gZsUEEv04h08xrmQZPXxe6IbjM2/gNw5ljz9/WMEHftERAc8P
u/75xHBOSx7j0FJ9j/FbpwXLTqYuyo9v0lJMg8arsb/MXGT2PT7Nby4ka79kJLVYIRx8pZwbIdqp
jjBhbk29rdc7g9nqKc6XiHfKdo1MpB7ZUAOIoJIJ9jG0QP7veOMi9YOxy4NQjK9eCc2uZw2qyf0m
36RGjttuV/NtmqKP9EacwdDJWU4QXZ1sxNiqlWamnaPEsDPcISEHdssHNRBzomxGX/KMs6ZOzvVT
xRYuLZQbdBRp52idBI6RdHwalMt3qaBqACwd6YesRZEHElZepAvzDT1/4Iant30QE7B/N912kb00
g6Byt8hbOkxF3UQX0mc7nVSPd1NsQx1LFRtn8KWnnpzFodvKs2PEEYX6H6q7gmqDQRxBifarIf0u
5hRCQgsYhfDJMD8vzw7bm4yXkltSxgJDAisAKtJiOccfNjUmMmej1tUjCVBqlL3MeFKrsfzT1PiW
NVXDiZlYcbTHFdkKxMD6jW6p8q6gvG381xTLJ84lbqv08uylMmCV3J7lk6ArPs878exrK+VOpawm
tE1BUc6R4Rhgfv6fDrhMoefDCxoc02izUm9Cwue9ELw0GfNShm0BF5AwIs30T6aCqLqPsM+bkSoZ
Rc88lzHJu3H+kDo8+4nmwR1GayEyUNPJWNgobov+Z9chQLjN0FyxG3e5vKRuPPGpxEB5JJYlIK9q
wcNv3u1bbM3264oEqEHO4M2RmNko0Y6RrLpWUsaLcTryVX4bssnFCVEOexmpukuLmizxQymXxqnx
SNTuFEb6UZYAwJ8AiOQeV5JWRMGbqAto7SxYRyvXxPLv5V43VRNuBiGL5SGsh0cHSv1HaSrDlhB1
YdtzFvtEKx3uWHWlyTZ1zPDfA/HCLSkW/EcEt95yZtNIG0f2/AH9IKOQ4F5ApYtQYCskTDU+bH38
+d1rHGwyAOomRFXT74735tC/y9y18RZOD/Iaxb3ZQRc1OICt5pU+k7DpwHszLf1lvTLaGlgdy7Kl
PAYMKbppUZRKwSwUi53C4Ay9LMhIyANOyd93a3W/U7syemfpFNmx1mKCFE+yZQy18DIoy+r9I7JF
YCbgh3+zzd/PRFgT986GKeUUHrUoP1yWXV2oE/iAiqieEA8u1BoSlgRaVrHQlHXPaiZEZwLxyMyK
M9vjtCDO6RWRa4t4BXt6Xnx/JFt6FTEz/bBS5DhKyfPlxra6UFIss6CYSalMnUOk1DfPgMYHdPx6
A/OS4g+3F/auPWiwddZAKuMXB5RnVaZyGVpqI4viOJAPGTsj8g5jMJejJDUKQCiqEV8SDnjgJWfv
qcJ3h/cCsmK/1o0W+k9bBBw5Ki2dzeiEi86ZyGFgdf5G9IdiRkpnqKZjDCcBRZXNSRboN5/bMEcY
jP1eiGzUoGjmDuErdEua7+fg6RFNPNn9Pn54wkfEGIi+YZB+81zG+Fb+zP5AgaW+VP8J3Wdh5sLG
eYdlw4o0UaimfkwQda/auflEfW7nIZLAs4aAXl3HXmELHan2qn6B0bE2lAeQLrAco8uZ5D0TqYAd
h2wZPLBLZa5CL85huLyuFldZVUiKmPm1TxJ7pKZKoCv1hVO3xGtirY939rLP6gElxGm8C2OPI+S8
EqaZ8ocWmcFpWntEguWYG6BwhgPDMh8Y9c8PGT1HRUBE41SyJk+IPVOIAwlymZxQuB4eht0V1mqs
Cp4X8o6wrHbK8PJ1RoMkq1xW1VNugcgFCxDL/HuDnNCK2mMcK+kcNSVNWlXshiJ7OdriCQ7/SYE5
h64KXSUh+ul/z1pfAUU82mWhJ9Drd6Bd02TeLcB3x+0AwGRH5sQsflqCwFzngxVs6FNhD/naVoWu
rRkL4/eqmZ+BXi7tuDCjZy2G+xmkTtFwU8e7FdGSeT5CAjgvU/lqFuuT3NAA1e00LW65ZZsAtyqz
TAw0+CL3iS3mEUPm2ae97WEamPF6AuAmhMq1KwzOooTw6CdIU4yg7wlzwNnjmCAFRYYaIFR6/vZa
jO4QRvL/SWICXgJD/y0UJw0+kWbupk+IUEfXmQeujk9jVTUrd5WeNbsrlM0IBWpMaTrIfFOGoSjB
N2wgG7GmgDSr6sWT2j/3s9Oj5AzLSEU76LOUZrVUQ1JvdFTRf9y7oQ7iH5bjeu91xz4sW6NGLMoJ
EZmFc54FWLhC5xXkPS7r0CQMZ1zoYS0u2Yi4vMMfvLpVRi+Xz2pBcU82H5x0KBtJ77UchbICMTxf
4UvzoQbxuxs3sdzgmlnDdN3ZSJOSgZVUn6+JRiRq+HEhuLuxJOcqgjk+buvkvGhCLDc33jrRWNaa
bMuaE0CafVPLegXVv9nUFToHjQxDWfaCNL14zi1HzblfjRE6pY2Ulfs6p16FsGtQBDGGgwFNob0p
PW0WmUDIHAcDAbmfCEpkdsDYbdryFkYGFPnN1F5GNfgpi0b5EV75qreggDKOaQcrPJYNbxQqaijO
D0LjTRLD5OloSE294DuTArsh2gCj4BjD8pMsA+TPQLwkOhkUkuSScu9fgPaLg3DLRfONC+SpI8aN
jLLjbUFCX0L3vhEo7YmwtKjRKtmcyS4kv+i7ErOEjNL9ss/LJ62D5MgYsVUUV3ebE6DqWj1cpUky
MFLiilUMvBZtmK9km20oGXTi/boOxw4+e0kjPgaBgpwRreV+WEBBU5EiwPRe1mJJoo/rZeuzFkKy
+3fev+HTkLUOdcULlpDuZyUzW6C1z4lU6iz+12u29Wil9eA88tTLltalVgsfNTLhiBLtIfP2zd4f
Woe5NcUnx+MY7HVXhpZ+g2a1jweDsLI6icSN190+q4OsC24M93XIhm+pieevkmM/lxYyuR9m52Cy
ebjAkzLbb4OyfhhJ/KK5DLWGsrqpaDF5z2LGqkRb4X4Ew7x176NVZLWqpP9Fza+X5sBGacz0fCbT
u416MvHkryCAotlY11xN3mzvnDz7BwsYemZkZzL84JxflXVphplV6CSxQqB0KZchovtdW+dzMFFI
N1y5y6icgYcqInaZmAZ1UhnInKuHeHgxxpG3OMmBQP2+Rqc3+6SjnTTUWYpythLlmBdz0Qx1S6B3
0HucLLwNTZ9s2IUC0OUheaU3iKnDE2XvVo0ycy2+Ix0NFhLvsSjyutCWipLWZe+LfKNQ2EqEOO9l
JG1J2f5jg6tDC7YFAbzBuJLTGdpxJ5zBr5IkAHWrAW/W2Mz+O11J9Uk54iEM5eccRLpj9PTqVLOC
8+zLgonK83r/gaMcifKwYLc6pHvKxbkAw8QnSrK+uIyzdc4Grv+lLss/xuvMe/dGZPQKJByfvgRC
/EhM1HDgQwWvEg2QsZnh8l3f+iahEHgO+Y4soyHK1VCuTz0RVjZFaPF2lKhyggihUJmzysxXkCyG
5HuXbVj2Ba6kYGDsmWvnQ6UgC+Kf5NBpbnoE7JztceUtLg+rA/S1FZ2chjplYi/yDgYrQObbmELd
48KFeyytjBLBQmwODCardTYBJUlSPboGCxarThVavTGNEXo8AL5W3Ko1QhX0h1F7y3DWkO91TLML
FchMI6+H2aZ0SalnWwW5fEcTroXAiz+cqvHC/kawm6/5zz7N4GUUhRpDvTJHUjUC1k/Ch1H0/yIZ
DVlwIQYeL+QQYrIPtKT4xzWeay6VFQF5u6AiN5CADwsJAd4wQt5u04kAimoiLmIfF5lEg49LMTuM
iPKjWU/J66rIuGtIx8uDswiueNe5r0UEhFI14rVQCpzWTZqsQ+rbxnZqaIzXago3CMciWHBbbm1m
KzSVeu9eNaIpQujjCnm2c0ZoarWh8rQRY2nsuxcZN+6rFYiJQV0g5PMnkdbUmMWQF7FMk6TlUyOb
mh6m03EVQqYtBTBjgBUO20YFVErMftFo8zxtWL6oYjJf9EmZ7HRXXacjewin+O7STj4BgTwh3RVd
8S0bxaBsHILoE0LzbvNR8KgURi5YkIbANuAX82YCRyheMlS0mL5dvy4kMycHp8CJPw0rW2/41b9M
LbHWH/Y1HIhEPt7ut2lCwmcfy+/oW4Rd+0BCfo9UIrkm+l/vK1Ftx0fnC26v1g3/cWwX4D02Y/A2
YsmWZWXb49Wpqcrd3O++DXLP1NQ4CNbmSu7wDfmDOchwMEUBCjytuKnxCwNIPSDlfSaayek9b09f
aV3gN8cbGV0QNM85xOLLFCRqLSXT3Yqs61+9TCbjO+XhWjSkaihSsfuYWwtDcLZV1IiYh8SUD9mu
gEQhqxrBE7iiAER3Rvrz3TZaa9WvFF0y/tQzSxcOmQjCC0bG+KEPeXiejpEOoMv89bVoGPvJ2IUP
4CJldzs9nw86+RCCr76vQJkiGlwofPvD0PECJdDonEZtt5HIUZPyav3ebLZHHKOpaIIkIo3bG5MQ
Ck+/gX6RnPZrWZvz6XynNdgvneWFNS6jsizsTYJR9u9hXDMnnwrpBsw/3RBH7EbFxd6ujEa0Umz+
1BogkjtjU3KT4GfjFYsDQl4KIhRDmu4ApUkPuPxQ7nfZs/5ihytzC0Tjk4VBA4YkwxOReASCx/hd
/0RCBjc/kFUisEjprtofq0UvOyFHOQerc2FH88MH8X8F/1iITRGcSEm1E3WWY+n5eZA/Pf0FLGpY
LL24yuN/iYOZstq/TLV8qv3Yiz2rrCoaE7LMg6MMYhZTnNmLeTxcxhVt85b76OVD07DZmyb+qYW9
yw5s5ea6juSQVaytWrI05CzPUEp1MCAO+G/eNhs/Z1nxWMmWw6jxNjmF5jawJsShb1u+Z6trvl7E
2u3Mcb5DeFdkc5V/kah8wZfuTk30VfBzCvoNvB16ebAYxuQAk93yg4pD1RS5vzGJX+ukLlB6vOkg
JBaB4T3325OpfMuSm7qTMMeM62YiVFTPqeL+76ei0t013/3grIWgSfX7qaAoeEAmBDvrS291Qu4a
SvgOd8yIDnZvrcMfCV2z40ZTHq3y7pO5oVRKuJaUi6krvr9ixPUCr/hxjPGytiEuG0/dvMgK5wSQ
quLTbyoob6qcGH+iY6eQksv4p/4t9KpBnyePaDgNHcJRBv01zqPGMvDbJHpKDIsGqcA2RF8cQb2a
TFlzUQXBOODl3c4HbkzOLoZN8dUjpFRShWu5CqI5j/B6LML6ldEIaKhIMzR6M1C5ibUH23urqo0T
Gfdr7rbXwlaTo+Zrgv/N2aES/kXEX/QBn8Fzir7AnXMxQ9SviG3aMuJrxioSl+yVy3q8RjlNzr+U
NMRiw6Ta0zXVE/v/NuDRVjj4b5xzf95d4n2pwWdYxvRB+otpOemjvjGh47LOQ9JWTr+utYTJiT5d
c0eShNxdNJKtsp0wWh7oqEhq07oViXlxHF7/02OWcLB+6PxdivdyTHrK5R2tSG9DxM5fP1LaKHj+
jiU5jZu7R8zkUXOkxztB2LG5j7uwbBLN8tK/mQAoYKaZD4j05i8qpBTfdhurCdAqoDIxm7R5JMk1
lsznmYpppUn90Sww0NJ5S0Dl230a3QjeuWN1TXP2IQZH7oo5yMYhKcAH5llBFGY8880Bdf2F2pTr
jfRn0KUGw3pZv43LboMps18vkWs0ps+hb7xOHEHYBJ7xOoCMtqToXX7Z94OU7QRd8kGC+pJ4simE
I6uNHKB6YG8tsSOiUu2LpIaZFkPe4vYHq/BWsh30KCrHveaBN2SL7+X3c6NKL5AXXRg6sm9cnoih
6xaXmD3aF+AEYTFGfn5EwzX+3UIXjXsvrhoM5lSGE4KBzqgdKcF5vILr7Z52PTFna2SlEjzSo1BI
A+xWpmvv2cGFivs699suYJ4be15W3cJ4ndO6+0nOarxkXsXM9y735saIyr5od/qUg6RnwgS1QIOJ
gIBTOrvk6yujQ3twvK65fFT5xFn8RwftQ3+uB93p2/p5NV2ICDP9RFd7gvHrVS97Gj/PzMEF4NZ7
gHRDUwAEihHo6iKjWn7YsKIgcMWVaV6irX9+2xdHJAf31QSBM53kpJXQybUu56wQnj4Z4MQ/MWyC
kVD7+V+hRemyG2kNfppT9gkCFftoe00LuFpxm6Wj9pExnd5Y2RWa0NrJbAyKohGC/N0UessNfxOy
+yTUqFRzmpJwIOJklIVgxHNDmoUhvIYkhK+xvt0domEo6hsKgUeWHkzme4MkfGMoLJJQB8SNpSol
MUFdnVpZFNcQbwtq5YwdBXxp2VnNan8LXJezoIeZjrVBuF+htAbyGUzcdW6MEosycmk+ua/iP+ow
vpaCsiazbt08AxshYWvrVvu+tlgRCvtIZkTi6y2IjgUxjz8Xh7lTRVOwzyg98JDWGBrttw/4Q4JE
5pYMemjcZKEEtnWS2cihmgF8ZzmO0XdOqGNvbDuj0URCS5c+wZT0+8sz093gtlI6QU1fePNRKDEo
Ayzr49KtG4FDo8+cA7vWqcIt5C/a1ZGkjSoGVdoMkHQ+OEWjHYGei4mdyErJQtQMIHvlAFDTlyL0
kOai47JH+JGU0xtuLO0qfEC4xjLuZaN4i1lqjC7v9D8xqy0xVMnDzFidWFjBQc3veAb9m79zg2Ph
bRmfCavuNXFajfGqpAMgtY7CRKAGVoKfmPvg2+x9+DordlOHE1L7VE7Skpz1XX4gDsbhhzGUZ8cE
D2vp6cMi9lk3gjjD8RKDygU2NkH2aHVXnnMTrLy6MhCtA1pL/Xo+qTY0jLhg8iK3O3vXfk59VNuL
yzCB3sXxJPiFe/gTIoqZHl2wlwU53eIKRH6L3PDUClaEDCfmtHvncOvCxQbmYHYLYHbeUDZBNhcb
3AbF37aD65gQqnVZA4/Scimvi5Hv7BOn0PMQ+zjF9nebXCqgOOlRC5+Nvtjvv3BHLUANGgp8UK2Z
aFRGyet3nVZ3CZVZtcKZP3xXQqZ3kqF0tyx2Gpw/XVrAotn8LsdC5udflD7yqJ89ubi4FAj5/ELl
va0KGEZZu/bEkGenQC1WqHfnHLVdA45+ohBIRaF2hBTzjYJLaONjWVmR12pO6MHKDny7b2ctDs1x
6ILu1UmMQBcK+Iz1vsKt/KKxHDUuoqR+6RdUy3P+0m/vZEHPL8rFK1GeSq/gTJ2Sq1Ibzbx+4OGS
yMu3sddgBdYjQiaFfiI6wKuwnJ6pj6vZ8NfEMAJiyS+fCA+QMf50BQLx71mAZfXpt6Gyj8A4TJ90
GRS7NTq3rghvcSIJCEg/Y4azW1YjtV8fEeXkFDD3uFWLfYuTD/0hjIZfqiPbYbstq7Eynan123Pr
HFOOwftsCzri49x2qAPpzr67lAp/npC0hvtbiiPpVdxb90JqXBTmbJUMTh7Q2QNxwn3h5ouo+EF8
qLPK/z0lHizrD7xrlpzwjPHz7eC085E1d1jwk6M6nRSuYJJu2aPgnQfWDlc2Q4OZs1dDB3Hc+svH
XE1uKsUKh6gSyXFnNIN4oj8k9QnR29WalNzptbKWxEhD8yz9Xq8E26m5ZqJWE4F7TA0uj0qNOzSi
1PjdG7FlLsZ9PccQ3Z3BWA5bZIVjemERYRCkDUfx4xX7GDJUU0W4uPxOXhhmzJmcUKnerXjlZE8R
u1SABsW6WENyHsR7NftfMyTIwQ+ddAnCSWUNMINFsokCDJXUvAu+9qWJJTExVWUkpwKDzpWZGMJa
7OXVBCxIiqUAG1nWHOKmzKWf5qghSKjrbpLlgSwDQkzcYT//B3uIkBsKKMe/LizYHw3Nznj7ymOv
LHpEPaHuAp6CeZ4pw/gv6/sC3dqa7/J5NcSnNskwzdtFKlmOh6hrMYD+VkcdbcqcUQZtBmSa3vkQ
tVTPe8jVlvWE7R8aUTDuj8E+g+gA/95NZD9/Ne3w9WWaC3N5RbPXHBJ3lpOXkuUP/Xx7iOpglLgG
q9y4erFCdzLnCgs1Ib9Y6oHsYuhZ3bWxlu9cPYepaw9HkqeOHurf0fGQxLZdFxyjET1hlsooH2SZ
ztuHEhWIC0HqXnk/7Tqfmbmg3HxA/QSqGST7ueiG//kol/sTj1In/EnFz5n6wdR8Mg8B7d6DLU3v
WoMSZ9CnIkH64S5emEzL1A5uuQVY4/pJQo/9C1VlS25v63EJw/vDTtuqGujEkW3MsIrBdMcmAIEk
g3wHpL/kwN/DFFAdbPwobH04s8S0lbaUtbIyP2aOjCsFAZ04h0Rb/+Lbouxzal9jI6d6Kxym5Z7K
znUhOTxzNx5e62uGupNcXKPCJ2giqPQIIX0UDdM3XESXmcZEU4QCr366EjH+gVI+8Hbwz0dGvnI7
fxSr7WPh04P70NNnshVTyOOc7sqhEu4jeWAe2asIZCvz1J6WNaG8aNrSV/hPyceG/C4at/D9W233
uG+1IyYwncLMxcmcG+Fgwb5EnFHYHVjHbBEV9pXOyuMfbbBEhGVyg0Msh1zvEhmjOmm/zko88Rhh
eV7kH3qIyMq0RRfQQ6ItM5D23yYYtPV4wHBxekj/ahzcL5FOKiO76fl9Z21g9RU3Tgnn8N52pSZX
QgmphCs1jJbt3cpJD4yXMkq3EDGWLKwhIwxfpjPcBdizGu70Tsr3YjpFN7cyh1HRCvUGNcSfyDbq
Jc6W6MhyKFHzFdxSp/YkeN48YcUHUfYZRS21Z411z5umE4mKV3tG06UzIcqqboRjgKoIu/X+7vKs
qOkN2FG+wQI2ShWOjdEZkBF4+ymrI/U/4OzKWcvDs9E2jq2QGO5sqb4qeh0ZeiMyiHgAqucXrc5B
O1hGoj3QBo1Kv1UkzOQz2ZXb0SCrff6DmqH9NBc93vRdxyNvoST9vvHaq0M8RC4Ib1luGWKGppqd
MpsLB0R6My29Ys4BwoFwmG2MBnxkkFO6Wj1KiPkdIrScCjBiMUCctSbRCa4VCV6npWP3uyCIzupk
iBZnvvt80d2iU9acjBRfMGDoE2di7Zx3Jr9Zp043BonIP36/PL2JJqV+kD0sEqE8Y6Wfy5aLrDWm
rGKAGaMHQHPdaEfObFPNjRyO3K4nR+IF/KIH9arbY1Q4ABzDaW7hRgxuTS+71JjpRtsIj5pAzDji
nVjNRHKgYkKD4yHGGZU8q+TsbdPr+zuYqf1Z8ReNu6yhKEx3fOs0r41mUerhtefwDvrYXKFOB6NP
QLRxZA6NPCMtMX39ZBFBpthZ3kXGRTB+rhp08PT5w36mahFSdMfq2tqMw0RUQn8Y1r8tgFk/wgSa
3sq/muAKFd0WCTUE4E3WvNQtzH6qDzkWKJXIBo6Xlw3FoBTHq4amRms9PdLkCiuTUCRdgPCl0eMl
sLwaH+E9lS4uJtIKmyUrZfyP5HwhKPh2/jDCVlj5FaYkhTFKKSKU6wpnVPDqZQWQ031v6pfuq39R
1JqvgOzV8gpF2epF8EZDNktw/dBbidplHkETQ5vWUK4PpFc+/0N3gHGH6hWRFpic+zNUqaR8AiUv
YWpIkXswXJ1YnQNc/SP2fWZ/oESR0F+m4wP7PobXEpyZ56LrF9+BD4bNDSFSzOVjM4pl/i3SEUVx
ZA8oj9gZP9+0L4D6KjsjE/e1xThauX/jBdF/e2Osx55J43xTF7cGHmyPayVtTryS/E6JtCYvQPrh
NCpqVo5RJvOa2WRHhieUKcSACr41OiOaBlMxc/21mLUSjhwtFaurO/j4fRhWzXJLfE+YMbcGdulX
bpi/BIrh86sSQ57UgM3EWw58FIZ6/Hd62j11wxlZtZHBmMc0fQtvMnMF9Yds42o+fq/oth55o2im
JTmfhnaQNSKh9N/gc404doYrkmdriVTrVGaAA4tFdzYEtaXOqqV4hcktXUcxw7pg0rtrQNxCM2cv
Brllk/qu2mCcqwlv1aFt/wE9tqlFOaxeIt7REVHIFUsgAP3ByKgvVr8ef9aJu9Q3ID1mebYQaqSR
7kKbdbevg3cIM+PHUJSVj+njpLAutaaIoAvNzBY5V1XANz2zVEgXkSf3JVm+P/v5cCLG5k5Fj1Y6
t1DE5OyP8aupYE6Xlqlh6pI3sNFRNRMf9gGoZ0jF/FnS6nmry5xwWf4aH8WqwVDLTNN1+VAjnzpN
Ju0aOQ7JypOIZHwIFP2UY2w0gfQbuRJbXaX+sgLcYElWvAnOoiDAPJ76/gPK0cHI0WsF0OEQR4Fg
O32b9Mq3J6GZfKv4MwSUhSda5d+FqnstB+vWWGh85wirZo0MVhd5jrTWXB1+5CLZujIlF/zOIAvA
CWGOKIK2M8CpGIc+UFrIN6lBCg6bp611CbCiTkALnJBVnuVUumuXbTazYF7EJLcj9Ax1yckZR7Ts
yvc9PSogVvu1aAIoqwhSXanMnzZz4Nyx6U7D6XHr8b3JCqhGEhYIXge8uP6pq42AZhwQlu1lJ246
4RWTSMMhz5S+ZQ2BahRQ+LODfXzJQx5Z1K4bOlAiQy+IbpV1GpFtKNqTgSjPuorGQGaHuWTyc1LC
gLosCPWFkky01ZyEfQVb3UJ601RU5E56rsPk/XclgXSx1y1S2rrSUjRDqofyI1+RyYWH0DuRtCBb
G4jlRmCBJTGgxOGhduMHg3FU5kNPlengz+FPpvgDEgWqK29RAblVGWKAEE9L1SIygSSPTSqoQV5e
ac4BA1Ukqw8IWWYVEEac4PZhuITGNgcmm6+SPPlvMeO+qmuuQkTFTkc89M4hCUbOw9eConMxS5T7
FBxpMx/htxQx3UemDySQbazSS1iEROsGn4qVqLUOQlpMfVqoB1JwZnDlVHrpO//xcDvJIuaOJmyU
hj23h3qhKeCDk/yCDDgtXmuaxzMfSVMowm7Q6V41gkkluq4B/lqtSw+47AIlWF4DyqcnISg2DKaQ
fvNSL013aW0iTCnjsppp7QcMG60DIQrZDX8QNRVHGEknnitv+QekVXUkF4r/SaHAw8dVvD4qL37O
2NxpkUIF+yw4oowraAWH2YYoxiRwNNGxm3Z3s/ZXQ0CDNb2T/R34k2xiwuEuhLarwecYb3bSYtfh
0pKM+D9q6CmlIy6AGqYEHYWGO04d3Kt22bkwczulSw6zpixG2pT0aAyWWfM0vqIe/i1eM+Oz8dHp
8sqH8hB/I8HmWpcigj9IzhktVbZpEFORfWtC+QDQo1GpuCA5wYzevKUDXLEf9qXmTEz4zgx7BZAL
aLkP1wiQSktiaP20Yu2H/P/72qv+xFZE4D7vk2gh7sepYkAYxqJ+iMArnYfSPHrrY24gV93NTUEZ
w3wLjY5GzW8mnACcJTpePKfuCoPR3AMnmJh/E5cEbIlxficWTGcXHwcGiVz6SQxVtf6Feisvyo8b
B9bb+yOBzffLIfbT0gRinGnaGLXlk0VAQ1VUzd6Y8m7bwMhYPdruZ4NUMih1XI6xUNtE/Lx3tS++
qqtUN29TIqy84wDlpimyj04O5uNzHU0yWD2Ng5rUp3sdNMc5HPBv/odtw+5p0p/F2DTC33EkGvgf
zm8kilrrtr6x+8c7RAglZlaa75o0TEVSivRq2jtSkvyCPt26gntZxwbizvfKXfSscAjWeIviovWn
11Yq7MiRYHMOaRJajkGL6zpXhPXaKaI3bP+xzIawnGXLC5Hxqc2Y6SAbfq/nYEUJByc4tRSq7sDk
AyqFZXl2XbTpQk4br/LRST9pIx05sLnmDj/pSi+nNP56nEonRWQso9GlLGG0ZPAFwT6hNutd7W+2
0nKc2dDP0XwynnKoqTGpioDLRI16ab6ipFdlTkO9DuTkbjE+DCv0BuiIRI+3WcOhe2qvcMBQ8CTt
TmjUHmYmumU2mZ2M7IrTG/3A4EQOopMCGM+36jsgeFHJti0HQU6sSViUkOtT2wFtqBXJZsgeBVY/
lmLIQyS0JxWkIUSePYBDMmRfUubAO55gc4rEl6Zhp5d2rEEdG1lqael7jm5Fgv3bV+Sm/jPDwulr
ZmnHH6QM9bzs7RLnGxZPVAKqANFlDeIR7m6IKYpgIKBgsIU9HeV9q2TUVHuuaK5vWquIvC+3NBAJ
rO23FEg06Hd5x6wpyVjVwWjJzwJgsqDQd+aoT2mCpPUBNXBmYS6b9Q3cCi1mOReDNtvW4sAsnOTX
n4LGLLmOTbRX3IUFap/9jNOuomUCMYsFvfcsTQvA8Efy1BgChoNfomXnYrBFEud2Rt01Fv3673YH
l8f8TIuhhaCnxry21vgSOIa0sViielz6bch6UIop4NWhZ4KUiBtYkNRWuBZshCtrhl6DMGTtOWez
G28w8nj+yqXHz/JHE8lg0Td4GNzQYkMuCJhddoGJbCz/I897m/FEdBrx9Z9+zbTveLxESc13fNU4
fjMgh7vyxmiK57RFwg6bGpzW3VD6letp788Zzs+7Ukuj3KY4PLtNi178HbPi0dWnw3Qo3ppdL1rE
jlf306hTI6MMgUjWSQ9tAEcj6BnZDj43QKobFYLkTpM/bW+JrGet4eY7onEyZ6/3SLIxlifRDu/m
tV/6BFuKliJtKgg0PMO1TY2LapTYLPhET/yC+JFwomAjWCbC+ZjFRyc7FKMm6LMPkkBRY/3ZuaDh
v8eGJm9uZ0aCWRvx9b+6ccEYqilMYJ+07Ba1mMy1f/v7nP7Xro8lle/UkIqAl2ET5x0HRdJnHyTo
1WCI/TOmeU97rZX9wcm0GVQ4jIVBWMWk5rQ0x4b1JNUQgYcjiGElutnSqa5LKIbbl0C5tyIjKn38
iEpym3n4r16nM378rDKyGw/93I55WQa0djNpWXs/z9JIBGzo9vhu3eJK2P/sOq6t90croweETmeN
hAOTk5Z/4Qjh84OKIMk1Su3nl3OgE/xsauURN+vZCp/qc+1nZ/uHL4gNLrcnXQ/makfBEgLKlWPt
GAMsdp/LSildtw03NxeqVvQfUhyknatjxuOLrly21E1/LzIIsuR0k+LApI61obA9kNzo2KoP87WA
MRTNkCxrchteeSHmnGrHjWxv0Kc81oXbJlkwaDEHXkQszZB9xBtv9MYtZMhCKFJl
`pragma protect end_protected
