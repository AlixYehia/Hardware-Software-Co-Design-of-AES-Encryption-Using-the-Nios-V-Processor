`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
NucjHrszQeK/eEFXbV04FrhPd/2+3ew7cm4pwP//zsv6+/ZL7m8LEjLmzWJH+/n/
hoMfHrQW1JLPYhfWcbzdR2C8scKEN/dn5pqO7HwJ43nmGCqJTl11HIvF5HO97ML7
UFOwy3NG/biKFUWjzMch+yksrw1DWc5iYmOEG6Aoljs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7856)
9cFyFNlYsKySj60WbvYkYUUumulcZst57C8o9+oaYO+0aYafQ452PGOuE0dRGq9r
Xrh5AFvUMPtULTvdzDKB2cKcafTdpjuqPZ8u+amzJJldsaGnAwDlcE7WqfXa5kBv
AoIeUIK4TMhsFlXD0PsGvBM8yEqivWvpLQAWFZBcMtmZP59+EiaSdPvlznPuxXkR
gWhCi4wtGfQFmrV7KHQZYxGJ5uUYHy823fEbb9ObvKwF7SsKk6uFeSXIzHqheWfu
Ob/nzLBPbD2gwipafwwkoqXHIVfd6ManPvaODtOE8HRZKJWUEL6VeSbRSPGAXEes
HwdOZMUYrP9u8Au4iqtGZ1tf4mio4gtM+rF7/zXWI2mmn5xn1lCF5TvNtcOwDNuu
qG6dbzswqSZ6qoqp7RNmEbdXbZtcqOa3AGV2rvAYdtqRlHcyScvz8lgY++UFdzE9
Qqj1b1DpF1sjGiLYZuEeMVLNkwaClYNibhfmeFRgtp2zABQ5VzjB91k9gKu4vdBh
ri6KmN5jvMlNSROFGGADHqlAOEoJNSPVlrj31xafXlHkE3I1S2o0i9Y1OtLascCj
vT+MKGU/L3Y5ZI75fu5kPZVMmCgM00n3yRTHX/S6RRNA9yiS107x333fZ7en5zo/
7fzIiTz7gSgGc2kh3LFzeZRaZz69cTdKkQnraPIjWFFkdx5XhSt+O2z9gV7YCOug
RJxMog9d/LSrY2SxeyhWCSeivVWG+Eivc7eIWIFQ5zsALkAG00OYfc8Yzej7RBP6
pqQckERD4Vq3lWQQVsZs06XyGIz7oeK8IQng010AmzIX5Pu1PhAwEpw1MDH5BKtg
fsGYPXSUKIkapkBlhcCfGRSlCxsilk2vJixahyCwgmFW07LcnUwbDjkU4HqldsKv
ZxFRtBFL78oZ3zBbATpz5QFB/po6nuwGGMABySsA+lcoNijDb6lIctjJbDSCCbU5
KWIK1syqka/xP9yQ3VnRL6A29i1B/z4eOjG5JQJOjIPpCXRNMgW+zr0elnkb5QSI
MvzCPNZ94ib52+Cu5BrM6wZVjyraG423kTVzeU00ac9v1AkaD6O+rb4NjrkqIChf
6kXHjQnj971YXv5TJBZ1CruksScFg9zR6ho/jIOqeVLypyY+3H767dqRNrLkgGgt
KgNQIVMakor1dygLf0ajF5YVPuM1gBYt4efCvgv7pMYXl6dQSNq6CE97iwWBDSKB
CYjXqsztRLV7q1HZb/+Qj1g5o9nl9JIMfIZvwRYMAIdYcTL60gcufwcEcBSEKAL3
ZzOjT3aBOIicHIEH3+xt9rQxM6vbLK7tsrT1dqbpgSQFcGYmvGFskxM/3SKEXhj4
dg+5NHbg/gr9pIRJJNnolzFBVXfLCRzFIUOPHyHXbTCsedhbX3rR+Rv8wvtdLPEA
WuDi4fYUcsl6FN3InTXSvFyd/QH+p3yLChhJ+42V3ogbpQ399qbno2cdNPXehMyG
OEIVU0wF20KzkAGdhkxMHN25ylIooxA7JO3Up43CxTkT++tatbKRrD9XnM1ij+QD
FmBhivWi8WcDBTkJMgmP4jdiQ1+TnfJJdc7fNlTxiNK8lAXZ0j2A91bEu06Qt4mw
kLnnFb+nplWy5QtuvTUwmYulc8yu0CY/A/osC1D23zNi15pHd328od7fDOb5fQwW
lPbUlVShXW4jCiXjFvuh5C8jYyd/MWXBQcveOzTVhTSZS+V6P6wxRjV2SDL0ccJw
NE7yHC8wsJJlROvVanLdVwWqOPoc43LkOped2C6T2P68VRIp+LmC4OdP8kO3fUrO
b+CO8DUVCniSz1XCA5S8eOUP5DNpfI7rojvjBEFdLddCIBJAO8Sr87wh9AlLicTd
MF4haKC7NJBN86l68TXWAFO6g0NnY1oLfKWEEsn8oOTPmOHVmyHld8TlE6ducAta
s6qYUaXqkoIJhf4YsBR4P5mxw409chEYT9+huFtgWCp/sRIKTipxeD84R0gZCXwx
Vsj4jy/UzLJKVwO+LEkLGrmKdnkh1CbmJQOIKNnOVw93ivjAUJ4TIN/IgAsvFFWQ
7xCJiFzXCnQfc54OEpiy7K5Zt+Q/S2Wq/MV3KkYcP7w6K+4/8zhFqAZoaqAFsD/g
Rm45TPAyRF9tmXtUbAuD/enkkL5m7TRENVCRKwTSGW/1liFniqEn0ny8uDlYl2aG
ihSGpGWAyyArA3xyjKw/v0ALqJ9k86af+BxAp9iRb/DF4x66CAvA8VTurrPt1G9e
qUKqupXLw4gxQmj3CsSdYQpKEyqbIdf+cuGRBl1zoKcGnDb1kVNHyWh1ncw1Jb08
qaGYBmwkUvlKZTJex3u42a4KTtqtmNmu+VzXKw8eJK2t+kAg49KEaZ8J9QKucbnD
wEJ8DzZKvH6So60h4p1peIUzaqFpegOr6aE8GLtxEd6H36HoD/8W0YXzbf82YZZm
wesxsCMu2iU7wLIJDE9JczvHk35PYSN+qIBRfuK440kHqF5dHwUAS3Txg+08aDuH
Swni7kgR0V1X6eL9vmv0ijaZ2Ohk5jtoOJK0vMj//qIUxqYzP0ruiST0TORCilB1
TCsTi5dIT0FD2pJo8KhsgIStNf01Jj1HW1ZpICtE1NAFuBsBYZ6v+XCBEBV2LN82
y/eZa92t5vs5wYjsN8P9MhuW1EBPkkLycLke1O6uOQKu3fwKUgrI9J7flExrVoQl
4nWswQ+ty+tn3LCIGbT5IgNlxedTvSf46A4TubtObjn339j8cnMxjF62g4bxbTAM
rcHSMpcTL6QweKiapVCcMYz2+yZmwyGRd8SZecQ7E93E4ZgSMwv2xYHn4OvBASnj
A2xSSLAeev1CDlS+wdCL3HvQRpvWzwK0JlhsTdWkejuFYfUwNkTCx3afLK2uX/Qz
sH7StU/lx211dpl0Le/MmAhE/k21F1JJ7iFiZ7Lr6viAlIvWbuCPaB1q+o69Uebx
+PyWGpiUs/o+ikWbyH8E8VltKaA8/xGDaGHKezXStvuYW9v3IwUqQemSOKu1AYPj
XcWSoyLLRK5VX+SafVzFmrT8CwRYqJyfXKUnC73GkX+/IYdjPse1iP2dPtZSfTr2
0qmjBLkb7hUoYAFyLXFWLovwW8LKI8ZCsqjMKDesPjjEYt44DmNuUjIgDU5ZoTR1
FQ6cNADvlCwS1K72ntwdymVVsS5R5ODeSRA+7krD73+lTeNzPYEmyl5Yzq0XjfLT
aH/Frj2hFRLcWabivkXYYZMnwr7Ki3wZGxM8v2OYxD9lnr+pP+22jD6Asy8YFBoy
txCU2tPMVo4YiGP5d2oy8Lq1dKiEObAPklt/tm7PcSBhK4KeBC0dlKit87BqYOBK
iJvu/NGYPhn4NCME80ZcIkkxN2W4phCTnfWEzyPxOF8TBKSfOd6eWD/mU6Ri3AH4
PxrybG//ur5qCaFxbh7VOfvjQDLYZWkI/1+Pfzpkc3T6V69RZ1HirQAArDRF1NyD
7ZYQNy7xgr7ZY+vmcqNybRs2VLhIG+zhD7IAk8EKFGd+oyEexdMtZw8HfRXZff1F
IBzYU/5y6YTjvt0bg9PYKhV6iLMZFecLEkEY8hlScjwrA14cIeTC84G5gjSWsDuS
GOIVYY7nkA/Eb+jfpy1cPOGhrd2JAsIqXFO55hdukVVvoNSxoKyYGUp+bupqKI7b
nkEYa9qU+mh2xJhAkzW7oSR0CmyGU8oDOuqom/nLZYpaBIFpFcNTgDqrf+/3oNuG
WbOiYJUWNNgsD6pQWsERkAkLRPVKm8c9V1akIxMJQ4ipt3BK8+yQH0Wx28PXXnpW
woGKT1frRQ/LXuXVxQS79jhHrlN08PZEG1bc0g6sGjCJXjy8OEmxilINMwpUR5RS
944gJp+EXPRVBPWumyvAra1G7WRIeXVi8wYu71TV5tF4w5S8fPu6qRIeFXv9YoHu
I+vNM264McDmbfiRtdmDV6Kj7/seeE4aB2lmJmI/7aDBwlYVE/JDUTSOFBjI0G09
jHcSTYM+mUz2fZqAR5Cm/v7tHQMJpsS8XsE5JoVDdPRcOyNiWFi+UtmFGaDlnkVl
zW+XEPwL2caQkTpf9yaNHplLeIOa36akpquhcntjwbXabxvlfxgshxWktwptG23l
TXvAgeMSH7kx94izwXQ0K9vIiSdtzr5t+j2pcmGRdJ/hWMSSHm3MpXNivTFlsynu
whJY5nLfB3tyGrr1XCfJhGjaY/ON9x9qjK4gDjEKaMlqFmLUgCF7NqhKLOnxS/Hq
KRFo6ougm0HO+NjmR02b3DTc0zTEkoJ17dONMBVCh7c2fQi6VlxvZclAG3ztvXj6
DLd6nnu4ydC7TkZbmSj8dV1gRKWT/OojojC+coPm1s3nrAFgRN2hSr7zsIaWG8ew
Lz3XD9QxZXgePjF+JeuDBjhZGioQGSIKApVYRhkvFTdB2AlBSf7D7Mo9RpYI9IRn
wWqdwio1cCbhhPd4RZB69J9/hl4INbcYP0/eLEyt8okbzrhguGuC5bIYWvHaOtN2
EonWBG9hexNppKYCInj95esEWXG0JyPKktcsrykcVEqBhv93UW40psdtUFC8IlHo
Dpfo1ekfTE8nbW2DPFRu9wiAqWmnit2FbBmkQIjld91Of8RtpyzIeCbnaQfb4eVd
Nz3ZwHYjQFtwRyX7Dn4yzgc5vSYf/syEgYtiM+ZuzJY53o6uxitOAOmOVDH9mFO7
9ygKVsCMKxEIY88+hhgTPNX7QdaCLeWlpvMQIKuATQXzCVEYu0qcbXR0n773O5Mc
d0YML5j290EmVAkLQ/7FREd1TknN26PqUEZqj1zJroA3KeYOnQHY3xnSCHlXsbL5
gT2T1XSKffRfzuIuBNAO0jxJT/Yd6j3WpBaUg0aZnW/WZketlVQObTBZNn9WNEDy
CUq+gsL0pdlE06TNKUX7jJmTByk5PgAuahI3R8ULcau6Xnz5wlfKhN5bzGvWU2R0
8kACffic0oN9tQXOkfSX3pyv9BkXZf3SOY7x6y8E1bRTBIqZznFoyqtQhxtLBr7u
fIRYnKGZCNThOaIfRA2jXaxjHc9wBbgyaD/1mD9aHNO40qeKDHiLDtmeU/qWGlf6
3E5+lW0nuLDLzUM5gXWTq8bb5py9DbxG3hdajFnS1TCPRPzVL0250YCzMGRTf/5j
9rPuG9JZSl6/bO94QTP2FOBDHn3Nq0Zy2bJpzomyGRqkKQ6mT2/1lT0Uff3ZX8iC
DOFsVK6afKDTeOKeygbscsPfIpUlpTzg5atz6d5cUrACVbLA4iVYVaVzEONF2HrX
yR7MSVUqsyEBOvVMXFK4arh7mF8b9SLIviLnuhihYlc3V50GL5+cQH87ZOVkRVmn
hfNV6/FM+qO/E46GpJGg1p39PoSSaJ8CpenBVF+t80Z5bZAjUgGohQw7Irn8GFn0
aeCDFXQT/zH2gP5mvhjdBoZ8ZfQUgaDhPNjBpEOp05zdfuStp+2f26xKL2kOSj9K
2/Jb8MFYPDtox90r9ypvrUEOxmBQsgtkZ76SbaWy++ttVMH6Ol4KLU3YP5kyio1W
cp4m54lOmB8qF3APbVYCyyWv7EiJrISwKFFvB60PNueP0GtA9ED3iSvw1WM0lq1Q
LUV0lZoNVzzWCRQ/eIG8tFfmg13I3yB+cuM4za84lsMV5ExpiZn9yBA6Afms3Cgd
kC3Dk8ixupz2c7WkzOFzIAHQ4AEt3lOhWeKsUrR7gLL/D2sFg+4nDC98LVLk3kVP
WFggNyXbF2GXYO4Mx8TXueZQjZo97PDMQ89tY9kTTOyB3WehrmI8KobHZrZna58d
74rOW6O2afFCedsbPCko4VTulofdXRsaWb3fkFSMiLW+GyEF9h+NY1KRqzBiufIL
JSoFPqY0etXfT6JoJkL8U7bF8hmv1/Yd3+5m6/QcdjdwFGIGm+dwxKx9TLMa0X3u
j13ilsqb3DC6WyX/mNE4zfM0ftIaeIwQ0Ed41n07RmSabi7JAFBegARRhtBWj88c
74K0t3WETmb1I4ukHAdHmlnrNXvd7rfelDZIjIlkGr9DuFHSQV0nK5IenTE6oPzX
OW2X7PB7OWEryLmy/juwnM7adC0qoz1vQheJC//LRPN4HrQ8ArUT+oJQzQJmjbeY
aLJ4FcsKn4pmabtjnnMc4q20805Ab51nj0RIYxQAeqxR5ubYm8aEJP0mAvZGMRd1
sj/JaDLNLwG1nJ/UuoFCc/fidu29eLqHD8pfUc5frhFmNYUAt+Olh8E03qmGt0Q6
mNwHQ/kx866/Tup0ejT22X/RQ4knvxNbJ9JyrRQfVd2BLnU66TpY/7xeJNGD2mRO
ZOlTAGpOeRKiu394GeROu7NYZflevecSdOGk4n3Db/PvFD7jUPZIeADpzu4nXU/n
7lQGgGNpeR+JOP0gq2BEt6OSOeaMBaW5l5IIH6wUP3f5VLToJ2Uak+A4CEejlMbo
4MpGiBWFVV8SVzTJofV2uqnLstaR42kf9BZdpqyTPqeycMEcXebMa92+Litx04Fb
/IyE7vHcfXIDbfODg0DiFTd5rJ7Q/PxzvwK87nvZfZtVhbOwREWQFepBd2ulDMJe
L5FL77v/Pl32dBy1r4gn5dcgfLZVSA0H6ckskxAaMcr/z/4w4hbLE/FUyAScBdjA
WreKZAwrDadHiIy0sj3PKFNs9omR6nUPW0tq7Y5jqkgVnEwgaOnBozSD9vT4dFBp
uZtBh0F3VPW0id3rGCdWAtV2/B8fqKMqwG/76HYGx3XoSg0f2zSZ+RAaPv6jqSbR
4gIehxPZXOF5R2K/0iyyvekK7wHaUaQwxnMcceEE6nBi6OCtJJvAZxWxWpB0KSXr
xkY7Q7k5tMloKrwtjKNl2fQPigx1xA9/JR+JfsEyfnyy6wY7wfvH3M93VTgaA0ZY
nTpMBRdBpacsbinhtkC323N+ektjvWeHk7NLAsXB80waZT00ocDI9+SDVxQkxd1b
w85SIgqFJ1KmRJoLZyzw/bOL+atZRRCRMTLaHEw1PMTXSMyMjnFaFBvjQI4kqGD5
wiwuV/QGUf/AcS2MVS2kO3m3xui50ezskMx2vLJhbnjmZ1P8soUgLwgRKqGjpId8
aYGjDj1XYbq79RCmqI3R8LAh7Y3zuGY41JhbGEMPqYpoY0M98xBxTjv/3tJQtruR
1DaacJYcOq/Iks7WX8u3SUB9yrJJr7+TH616wk5/8XEu7gYnzqh+tUkL6yjoqH2K
MCJt/EmiKq0Lp7Uoh1mJxKi6N9m6KyEQazy1NSF+14bQEhVFaseqHGXjwsx3UEdE
jGPr+T8YQwafTl1SputKNr/lu8f8ZU6k19FBHaiFXxNp2AzHeS2Z/lvCQjamGRsf
HBzWbVHo38vALe7VwCtzD90a57wJbYdi4Vabaap+hJ9Sul61ghpQTg7xrLy6HZr9
TUuHNxFFDOceb1Qy7Sboh1u8836zoF9CYdgSDu7X2M+yhSgICvrt93KG1idrrLx2
qkFm29cAvHoUQog2gLiwIfumgEpnCRP7boYBX5SXLMFErq+fDnZ0Wf2ogY513CXX
DgJ1whL4XFrEw5YN+wkwoOMCsIbOxjIzqwGb3dTXP6uuWUO2lWcWesM9Ev4MHZp4
obtbKqpY+rzYsfyYT79bobWpefCHns3FeRNirK0VxT6pIIbsFWDmxVH9I1k8EFyX
Ff+DBw4rNFyv+CU6It4Dx1W8m8BRtjpfHeIb9qv+KWZICMAVmcDn4Fxqcm300VX0
LXDnQ48QvPvT3ovWNkQLM8SvBa7S5lUoj4hLWByjuMfxdgO0asJ2jLa8UMq9Iik4
9u7TSq14mXE4nVQy6fvGwQBzG/SW2lDYfxF4ogr2QZvoh0PvCDW+Pe9KncyBXpYv
mO0ysJ2FDBb1QdA0HPkiKix8jj4tGNhHFvX3HZqdKYUTKKYQ7g01jhLmb52u3wLP
9pGU2WCVVT+9iM4FMiHucTZF4zJTGukmDDISCXJoAhIyu8s3yK1qJV+B0jk1uUPD
zs5irpDCQ4syHKHQMgnRAm/5WTXq5Gexdo+7t1BTfmvkXWiNSIoihlwn076/qpWV
WzNZWRwd8t8UtirHx1DFaNync2NO8mIWjJUO6Tnqd5li86BZUutlCC8b5nZEWkkq
pnbFEaLFY1EG1tZbeQ324KciqYtZzYwjohx1NYkB58W825vaE0D7qHK1xVi0afMU
5RXe0YLJt1+ZIXR2neUG9U9z8oiQelGQqwdA7cVaP5LdbLYavc5yxcEYTy0ZCzGp
hEz5Q+HktGh0v0JPBpqUhA8/FuoF4vKhkcSkNKqDHZ3UwzchyVFqW5LTQp7hFhnE
YGfmvaGPajBVf+stC2+tXBdeVvnP2rOGnW02GX2vD/E7gjX2x4R4U9X9MIt/d9TY
Oh4J3755jm1p7hddqq+4YCvJ+IYBFULAhkrUa7PK3TNiadnl2pPlVJhWX7IK2ynP
o7ndJQwV7CT4OM16A5u4Eq3u6hqMyDA69O5VeQ4fKVacKzzTCuMe+9IyIUWGkTWf
81DDi4Po+JuwL7n2DBzxvgX1jYACNO4lXgQj/HMpS2yn1ebEAdBs6NIzNv8DZEDN
N4h0FSGmioYInd+ViOIVxEoMUeSzgYoCc1UWzaT1uhev0DYugrV/CfSbE830EB9C
upf9TaXcUx/lf159ZHipw5l4j9Dmuk9U0ROqxQgX4MrYbjOxZuBMnOYQGbf5bElz
N/Emjyn25voP/cxzN9nPTPSXXxKOwncekaoD6Av4KS93jtPflqkV+/Yf7HIfQT1I
SWJ8uVRFJBXMxtqBa8h2hPD486Hx0QHx+g6IzocgpXKlNimAV7GH6pf59P6s/zRO
/NEhJWKbykVDoXrZPpH75LTmVVXeZ36Gk2dCxaosButeMH/vSi4Vj+jjSN3RDZhD
EfClqB93zw8/3vck3KjBA2iHQpYWiuT/3qdLg/z55v2E8HW5smOw3+YJ6xxoDHtB
J4vWhGgI9I+OdIN8YJFnQY6vZP+W/++P+nczN7t/OLenmudGCxMCmEt/23gXgTZj
v0T6VZtvaMkbkqG6WI1MnaudBQPXsT987tUOuXmBDXMfUYT4JPl1wgNDosSjBsIh
0kFxyycNxpYJD6719GHBXGua2RHkeeJa4zDz+WpYUituxF17UgbvvoFvZ3vZTE3S
YuuJRsFyxd/5RFTHxuArCFgQUzshUxtudNN0JuV4hC6S029Xf+LQ2kKP2LvM1+Do
K8MDChqgd/pRMLPX2NvNZIVHctAAtZj9tDkKYTFJ6BtPa1/UKH8QZefAdavtwA98
cwcuub5Tqit5ZsBGQJVI4Vh/9XPkTns2vKxv56shymWt7w+nD6kbUXZr+tf4tn+N
S5BkfMXd/x3NDS9GTTffk3psvVKqvUN6s/Kst60/h4uUytgCuVvFyrvQznpY16Bq
jZiDo8VzN1nyGjrAbJeQTU4ePmknfYxt1Ne161v0mBml5jzMwS8OoTFtiAkbSwKt
1djq+bvHPqba5A90tCGy+jX8ipBBPJOfqWFI3sUFVxTTILNSspLYoiNL0JmVBw4W
Brb2StHuqxyml06Mxh7M4QqfibhTV4rjHg+YLdEKNUB4OYLIqop06OMY6xSbGcqC
Iqi1naG8gE4e4CTbo/Mpi7R0f0eX38s/6QIgZgNtxnnQXn2IvERkzTs2+H5x6U+o
cnxzNXwRe6mM/b5U0drxxHizwzMtnUwZGrbefb9vwe2HNe59tAWWh2OQZX54s137
Oq6d2BqnFiKqgOKeU/sOUSo1l20FBjIU7zKRAPynRP+pAahgOSSi0PbYhcH7O/Jy
Na3cjYJrIX7kCjaQVpd7Egpd/qV2BUC926fFnOb6ZPSPTBkCUk5ke3+wU3UpxXLv
IzV9OGrr/Hyoh0wAdPhFO0hIKFPK0q+C8G7am6JvsMjaMSt9soZ3aElbeOdvDkIH
UiRTl4A+H31usJ8TOPwyAt+AWMHBV8mqSmbcgB4IGorH1S60O5YV4s90jUL5GmZ0
HQ9Buw74SxZAiTRX6vfeih+75qpsSrK1cJ9KG+WKh2vb0W4LIgJNjheqfjIx+If6
lk8MEkAZfjx6n3KFuFayuUC7ollUwg/JRn/otq02+pOT4fvHLMhvWaNvuHUTdV+Y
7pcTH+knTQqQL1mSgLdnpnuI7dKB6R0KYWOYGWoaPeh46NVONLRxoECzfm9FDO6G
aoNhHvMVd/VlnKOcL9to0hTrgONH06XJATK/gBVXMVtoef6iHkq9PcZWeH320OoB
S41wzte6n4vD/WbDhnBs/on25TsKfmR/uBrXTcTxxq0RbvilmT3N9Dj6Y+bNGXRV
4u86iWNguCotGMg+ynUZ5IryvdMNKnVDKyXtKLGMysOxnVJaBCaEQydy5W5CpN5q
VqR6jGwZfXYIa9cbUytjJYGkNiFCqZ+LmkyMFo6c4c6DpC9W2dZtRoCc/zekrKeQ
+zMRpeANYbGqTtWSs0lrJCKF8nOXsh2JhBIrNNteElhEa0L10sMf+H5j4QI6u7OG
sjjmnFYOMuZDoJewbWDjhIyAhq3YJF85cydmPS4V0/U=
`pragma protect end_protected
