`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lMppebih1qsMn5Pt60YSncX3E7J9MgRtt7eBFLvwxzHbmZvHTGBC9ndrClgXpHET
BxRwwhB2w1vTRswrlMJRiyNnZxyQHcebi+FMfFa2quzs2mpwTYRuDZNm5n029mqG
IDrbgAe6IgdEQsPRfxYm1pTpgEfrOYUt59UqHHa835s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7808)
nam3PRsKEFznt2gyQSZwKfbzAp1TduGRhAX5vSfA77n2LbQiYyMEBA+j9bwo0+oA
+FDB0dETXKFNdQ+HvJaseEbWhF8SIYyslLq/HLNerXEUuRLnGqUbRQbzZKbG6ePt
JEDbIymEHfN5lemZ3p7nxjWiaSJwx/TYvisLxcDg40X5Sx2dfTJqUooaTYynJ5z7
ac5wjbVNwOmoF3PLcJf/ERWHpV4yEg8j3E7AZrrlJk8+cf6LeIUeL04nPUqGWsyW
nwIU0xDEzvAC1Jtzfv2MB/E9oLhSdPPNv77Q1JOm4fNdMR6X054/KI5eRIqgV9Mj
RiAwikeT2IKX6koRYmtUFNNY7AbdcgLh5JV0RadUSucTemrU0ZSuPqXF47yjhLTn
1vO7JcauuUQw7HvYObjesP3+G7inM5k8vsqQCw6dw0mGLhqZLOBFz1P9BiuCjP3w
tqAJfPUtebp+ylTD9xMeMUA789eMGfIOsoRaLlKQAp9IZ2Y/LIvFke/tPVa7sTY9
x5MnZ2ZVxIXW1Y3cRfBYCWKVy/y6vcl7/BYuDQgoot28b6Qy+s6nz02MdAhCYe2O
xf4upIs0nLJq/cX75E57rOfnho7yM1g+jsA6SIwY2g6AxIrqzB7u+K/FmBPmW5Y0
jCpuvS3D3qZCay8qMSYAYbrmjvctvYxYdAoyBP219H0qUvtIhoiosAQQykYR4nZ7
DETQHbzvTSbNcHNBIPqeNBQrLy6wDK53cDue298ZmbZFoVNPHE3Lzbc+44u5kP0n
AMunOulBlFFNevF3avxZorKa9zxPGQuzLjbrPllvDYh1yBKtoN+oZ922MmPoT/v3
b+q0Hd5J/39oPLREUSNZrzTKh2xcZ5mRricpSQ0fN2SE6ZcLJCkDccbqEBy0XY64
foYi319Oc3Rk+3dmG8weUeD6E3aETAiX2ALzTj0AlNrNFBOcFhq2rDJ/ZvudMBgd
6SKH4ynPFfT/B6cg+EJFd4a5/nW+lCBCn0tCnp9wseoo4CyIlevpGU04qS3Z0dQn
JpP16vj83NLDpPrmaKLCMKrngXffkqYhhauVODJTL9/LlgqyWNsF1hxYqyabske2
oYkXinVc/eo3CKzSysi0eBuZbhGVeG2dizzH3zGe9wI8zGVjoqW9rT9duBOrXzHK
97X+o1ESBhFU8zyCLvYXA+xlxd2ZMbt4eY1vR6mv62YShqiJK8ZOF1m5oWuxNPqk
4jJbX+Q35FEzReOmCLZIW7uxwEy3pjgT0HwgzrpVh18tdFyqgs+Wz4TOGVfEYXqH
12J9wHBKtqIo7yZdJCQliWemHoM1P7lPstCjrgD6XptH6yYpkCrq+BEH18xwQLZJ
CZ9O7SL7E0TKc2NdEV813Pcm+vQo0fSdDmfHlAiOi0nKN1+Erz2+nyTuxWyKotc8
azIVx6rOndWBaPzpRfaCyjrvzq4yCYNCZyoQob6H+Qeb3tKE1aMQ4S2ypYfQ8CNs
OlfiPckehU9rSj8cG+8waNIhFU3lXktO1YNH/pETLtBQ4zW8s2vxmIJIjBhycLuo
CzHnQWp5DsTh5z19bLLXQL06L0nxQAkBXnYu7cZp0HLyp9HZWl319/17pMottKXZ
HjmIO172Hg2+7T6WmxhSYm0ih9i7zXE/aYRY+/W7qCH0CbYMGMbAcGRT59ktrS8v
9O2RJtw6HfgbqavdWNRJRqLEVNHFMk/aAWCzmRl7XuoUicTkvRAUCtv1y1SGpfoI
SS0C8TxHzSR3umoZLk4nOL6c/+HR3M8VBeXFuy7HLUZ3IueTPceY4Vnw3gtsk9qa
/wgPy3PozRL2D9Kb1DOWa7qnfckpIpSvDMMHRc7ipHufaAue7j5hUFLo7LqZmwWw
wU9tt934RN4gF97k6cawCrGqOo85WnMAgVtbtGpj58VG1WGZ0bwaIHL+FMHVaZHY
cWTwEHVgnic5aJMWCdsa11WkciNyEjBtbkL/78ZYuRUWA+os6/iUk75/E6ZWclaN
5Khs90Nhca1jE+DEyMo2WCR9wKIYrKoJs7kK9k6J8cEPijBwD6MVWLGDGeTLMssU
Y4iuWGdx1Xn7KWJ76N5Uh9twwfcAvSLR3CE5ptqeXaqo410WxcY3ko9Z0mP+sgmt
mEBTY9xVvd/fbUGkPvwRPRxSkLDwn7OFQc4ShwlyABZHAgCLGMgY9tdtyXezmnJu
nZ2tnoaFLLk8C2uwmbZWrBloSF1AbzrP/OSa3L6OruybBJDvot3P+3L9fsxjBmqg
9mO8qEUtoHlvuR7F7r9NgtapXht9BAoPnHqaHiOCiFNV1hXQAucqXHPV+YUc+LPa
Ze13cqoRAZ2LzsevmbYNxYDMH0TlyoJpZcZOdJwHK796tJifesFzbo8i+qqlm0N7
y1SCnxEvYEcIm0P8zWapOYqDaGnCXbC/yODsiSkSfnv7oQRSy36KnZYVbRJrhZgx
IfWxQ5TtqClKom5to7jUZVztsEbPTccWcJUXmQGrGRX3fnyF7+3aAXjaEXzxn9gi
aZpPh+MLtWB6kuqK1iqWxkiCyFh4f1VxuHzE7c9EJPtsV9e/aBFKwy9ykJlXyRgQ
KAidZlepDm+Eym872qPG36qKw/gwdjjYlxRZl7jwJ+DZY4qnSIZVC0O/Q6WinINC
K9iwIf4df00oh1XyHtTlUBJwDjR17YtyjSmQ6CyeDHo47J28w8sgut3nQ2h4RmCZ
tZq/Wl5+enjRwGn54UehXNoMhVYZkehtV9wFy9HiNrC1KjWiWOR68o+KLW4mozY8
gt6gslksZK/P+eqnNF1UkKyU60+zxNe365FWDfeH7dgteWRnIhuOuorxqlQkRSbn
kHBVdXgfTDjdZDKDXyq9pbU8ciS0CntAzXeMjDsa2QTHNVSKG+CcGfIL6VNNtq/t
PcKOgLYqB6+zNOsLjoL+j+2diZDZJ7OaYLb3Z4l3bzINSI7vh9bDoA8OAthak0Qe
ICYeUuKfq62YpDMYzPUi7iAplLnGKadNNUj24TV7KwAUCniEO+kJtHGkclQQxS+Y
3xS5arQHwBDao0jvc1Njg7LFt9fp+xyPiN7elF0c2aoD3bYqefzkg6HIJNJYb3uU
d3/AuPw+vvut+Zki8hG90jmQjkCUmUj6rqa4FeAbwtOu6oXCmLLutV9z0RaKOKrz
hUQoCQ8p6FqZ7QVqLWQ5esmhm3dNX+91OFUZo8dgTQAirY2hy6hOSVT3KS5SSKuo
PyUyv1QKTQxvmbBO1YMt9ntGNH29bLIzblg0OogaPR0rdpHmV485Sr3sY0twHZXS
V5+58dd+PS5YVHFv7DFaqSxF72HIQSyk2UQmboukoBWhC2fC/ipxwlM7C4j3e34c
ZsYhe1Im+UwnxKUAQS65uXUOGAFXcqrAH4taNnboVy3nXWUm2hdeTv2VPHGGIsFk
KWmWbC2XnquZU/IbZWWEQnRJHybp+jb6joX9U5Ee2xQoUUfZYOscCssguXdYRILo
Munc/f+1YDVckk6O4c643v/vhEjrugnJR5E7/dqo91dvs1dqzPHOp8CQANgNhLv0
MvN6i8X4ZE67c+lwsPOTWYPW9AvuxC14Wn0pXf8p/BpFKLNOqIqWBcgtUweyedDb
fkqGU+MqSGv/tPDlnTOTc7m3DL7C0N/3U4u4DU+ZaOst/765kQqVM1DAuKktsMjA
HYhzuOREpkSZ2/mel0lpFXNbTQr3HgjfZwopVmcF9yeH2gRx6pAhgvJV2gmiPfew
jxEG1KZXVqOzpjfht98I4hp8TLq7PuGXtLqPQ81ZU4p/GXg3guOXzP07v3fgIuwr
M9X0BrVCUIhv6aY6jWhDMfXvm2dmJgERXXbZn9dvImWkW7GMoKobRTJzjRnNp8pS
9xGjuo/CcT01YZLKbNjRC897T7kEaL5u1zw2Kj4dqvTAMEVHVEctHKVYDNKlu5EG
+9FKNoE0GEgkHPIKOtejfpb28Wz7fc+dDNRlDD/YIaH6/Sl+ZV15IyWW+ichgOeo
864RJFYrgjbEw1QwBu+vgiRelacmflIK3rxUlkarib4F65s18zKI7suoMriLCqRz
f7nMJ+hJ0vQ98Q/4MhbAdtDfGKdM9OXa1BaBY16WZcbtRcJf2ypoTNRp9GY1oC1J
E7fh7x/TiNf76P7V4f7ftTO/YWKut8NoIV0omJePFLJXlSTIfdg1459HRyCZCVRc
WsfXH+3Hj66Gh/P9NvUzihAo3Eh7iMoXyMOg/pDpPlBiHNBEPcLIJRz5O6OERUJT
vqO/enx3be6Fhf4nJp1NKxtEWoKKOEfrEAvVjmUGdWXF9Y44COxxDsH44kJDRoNG
vud4Z1oRflSXUQlDgM9IzrCn6h4zdwumF8foLuZjinZ7vuC7TRbGB0t4lFHcO5dl
leKdlstKYomG6n8WPsiLtfhtXHd3PB07QT4tfza36ufGADSuQvNBloDawH79Kkmm
ureueOrqTsnmyBuc+XWegV482v5CE4aSx2ae834zATwYWw25ZzuEKU3LaV2z5WXb
PpcyY8Us6skY/1/QizdvYvV4JoxVOaMhbkjz2fTstic1Ci2m8kKRZlwlgMy3bQo8
12yjCjapCKkMT7/KJ3wSEPI6YwDuBOo5T7usagyTFqHNAp2G9HYMl33wia3MRzNO
RZYFA6iJlsC9vhKLdQ6Q6fPLdCBn4s77uvcP5UFrZpqs7a1GwsPQblMt/Y3UtOO7
/vFLLFXsBI8e77HAYFVh2TGJGS0EKSi0lqpEMGqGmnr5AnP87fzW/y39NExUJe7Z
IbI+lN9Wa7nNHoowFrla0vOXEmfvpwR5IFyTQVr0I1ZmoizIYquqLSsjGZWDN8pB
wlmthUa+OPcUWdKNTZxZexLc/enTJ56L+tvXF53dSMuN63afsz6n8lxY2sfVjHrO
uIoJ1JnSIvHDAxpbrd8fcAUHsLq0DkN80+WQB6ESm/WxGKCSPWawjleqd3/81Li7
pIN9rpHM5jk99dOmIvu6s6pXVnrBktVStSQ5SA4wErVHXz3MXdmb1+puGfYyQQmS
jkMkanS1aqPOt4ttN3g0l1EhN6F7JGnR0MjbVbhV/ThdDCuK68cqJ7sK102vq4kM
AhBPGH2hnNpPL5Vksh/XUUaWOP4cXOxm9BWai31y09cKcJ813bc/vQsMAJYgmjGg
kachDUEBgYsia6JHTfT2r8KOyfn18eS24Q1M4ShRqnM7PN6CwD9iw9QutLQijVqE
zRrkM2CpBRFN+YI+AQJno8YZeYFgUfrtc1ItKmJOiSGhT4+eiGdohEdDfc8RjXwW
yieMcE2RYt67UIswhw8Ilp/67NCLG5u0BKMvJIh9Fj/erNG1CKiIGjnWziHR7win
BjVLZIGweHAJ6sba7sOJz/DjMXHr7yah8k2zHVBQlYfx6F+JYpHdbsdicW3wV6es
z375MPTBl+L5DfEHJGuCTFr4x8uNzi1EP9vt8LNQj8hLKGaniiOhle9pPhT8Yhfa
LuDwurAm+Aba0uefuXyhnz1Y+zn7ugteq6nUMSHVYstVI8JRQanQYD6iVPJOl9m9
43GDHnELfNDslTDQGOcLrOTVXxjsSn9EAC61VD2UdUy2A/b27Q9UTq7CJLTthGGR
GgaA+2VGYibuFubiY+WOm1F2uvXWVmMWecCo1W2/qW4S36Wgp1l54VCLyTbS0jfb
cg1pgPbehZtHfnbYVTHZ/292nusE2gyHHj3y7ckXpZ90LdokVekQeMs/5xDBMd34
OyBNvOC4p853PxVl1oCYsMWPK7+1b2VxL1IWzwCkKTCxwd6LwGzNcoIhV9X+lZgB
fdvIAakneCsxZ8pC7fApWBsUWgeudJ5ZNMRT8AEI2Zdz6jb3aoABAKKYVvP6LcID
8ZXi8aRgmqHwJ6L4vBecW2kFHNKEsKiv+e/vq0AjUC/XQVwscJdRZ5VcNScsn01g
MhpsDaPR5UPTHiQN4XNjcMbOb2jSGj01zqAoMY9y3JCwdrUP8RrK9lI7CILKMmYc
6ZsoNIQXyxoEwC0G2OrXLgI4hv66mVuZHo3RMP4F9i4hsqyYQSiJs5bigKc9jOF1
pPL2Q5PIVAybLX0JyHVooio+WKGZvDUDPeJSxHEHAlbofp0uvfzWPV8e3E0t3fOY
e4FxIdGFLoYhbzhcouDR5KRXqdo/FXOo8yoeun1JbnA22zxX890jMj66n8f8ILXV
NyZWSgCmgo4FMKoq5RJ3J+eebNfNIrbKtlnc2r7iRbFHWFhWanspjogzk8NIqUDt
gmB0Tqhg4j6CSPYBW8iIOHKt7fCIibiJjIzcDWMOPzJRVp/KDwEkJgQJ9+u580aZ
9YST5LahkGB0FgKddInjQ20QZMgI0z5o5n3LTkyiBb8eCs9I7P751H6oGcCPuszY
iYs43WiZA4n6mgyIn7fM/bJCCQKrRuoU4uEvTAiwEwPf6tuDdy6dD9V+ByisVV/n
cAo6PkXAb1hCfZpEU/ybsZwdgqyZR0NKWleIEsqST0C4cC3y8xzMJnqy5rnKDI5a
u25Qi8+WNl3sb0kgMcTtic9K+X1CaoSZN9XMXf+gLGjNSx6YnYii0+JDmsBh7prt
O/cvK19HvOpizE90ZPCNoPY3jPDWuT+GCkp1ADC9yl1FIvFyq3Zs3QQnvJd5mgGn
439nebo/eIq6KY6DZiKPzCFiaS4uhCB9342/F4wo+8X37mRlRdEqRncIDuc1Mrvs
juGUWvkQP2t1634O8bm9GKFpCe9/1hQzS8oNnkiM1e46kJ/vtN0rp+JnGoxmtEkI
esdgUz2BomCDmgaJasdLltSGoKg1OoRokt5Ct7p/EBOKdVr/o2Q6agqvgHq8TEKy
q4LvjET4xd3d4sH5XySn3wg8KpTtFW4zSYrz1kWq90S+6IJHdNTziOJEcb+761K7
nmFqf+xY/ZrAb2BOAmTVAm2ERNH9pt4c2bPeCP6RF48O6IJ1A3DDirxR6FhAwYVY
y2C2/ftn/4NEKq7knFaT1fKsI/h60Rx+B/u6DZARMfbjA3rfBTtR8E5pPkfi7AsT
53BTMPAJGnE0xD2sVGU0Jen0r4yyZkUp6dtbARyEAiXtM/2aZaaNcup13+2ta4Yx
cCh3amc554GEg17JPKd/6bv+KwkUNqGVpxtjtxZeUi4ttE4xyJ1py85PEtoosOwv
W3kLhISmE+8ljbrFq1Vr8YyQVzVUGzaId0yu4iGnqQ6Z84qDsyI/gQ31fvTiLJuG
twx0JlGs0ut3TQoua0KiQsYBrgy/wPOZ4yvNtqeYrFt9GjqZdB2e6W22znpBZRqh
XhzIsisEc24fJvg7PNIglnkVUaIOVaYnQb8ZNn7I81576RgvC5j/XbF9MIimHFTY
TPf0lNe0w5Wun3zqRaYNDj6n7phH0orqf7U0NLjhVl4fwCuwErZ+ygVFHp7Bdr6l
T/k3vhMdxSYeTIRgte/kBfsX5TI0QPXbgmcjB3b/VTG59RijifQEVSZoCVUun/I9
aCkN5AjjlltMLL05DEF//GQyMa46i9UbEM1FstAohsiJSuHLCbv9Q9F1p4dRDmXc
YlY0JM/iKOtfSWglcCdloXRrZqmxJgsfmygLTnd1QWk9VJBNfgOsYld3De5IWCGI
cRRuiyjnRm9qGntNNIyY2M+tp5I8Mz3kuSJBiErFvAOACJKhpU0ec1dhzTjCwWi4
1BZ5WeSmL/A8ygCByevNiVqMq5xhE8ZsEp7ofmoF05LPb+LwnbNP5Z1xmhcYN0t8
mVbIxhkjeoLmhcGiu8awrcxAgHESBy2jbK83H898/nvRPvhR3jOptiuMdzBjWs8r
77OWRT91RDHAs/LvrWrBjotPslin3XbaCEGzrnNzhWMt19l4K+ogiUz00RVGy3/n
N6bkRK1jg5z/zJ4WaJO/g0iWCZNI8G5fASt19GhopvJc3Qi6dDenLYHObSDUnprp
sx8wf3Fmjx2sFp2doYNqmwGqKXMlQfwb7FKO4G0HLyouM9RGHHuUTxQvnu1XnmEP
9YFmDhxRRXw4nV8ZbDzHSjQ+Ecpx7bMhtNWq1Szqp95FuCJsxENilBt/hTaBZ+72
92B1OQngHxhpNyV7o9sbFwN8d1RFGy5BEEURwNb2NvJnqmFmXuUYRmp8Zj+L59oV
H0SElxlH5SbLWewwWnZ6WCh/6eZxCQtoSNy2KLrC881omwZsnQqJf60Loo9L1OoY
37scCqJ6BjkpD8vry1Wnjb7oGGPGoJCM4UZvgmoAH4YwPqC3sNxb41HX9OZrBAM+
pbST5/AWtTH7YySs6qXM15F77RUUFImHczdNL0bDgCfIaccjb+i93zM+bzGmzgWe
lMnrec3e6/wUR3/Pj9vhlyB0H1Mwc8/Wx/u+iGjKZVOcEbwZPGBZWXbjpQm3rDce
u8+kxTdzVSdRi1tRI19g8seYuRz4AWZBz+bGKG0sWdfFf0ru+seCzh4awVM1XprQ
RoUkxaeUKGswqNF1zt5oPU6+glITVNzh9FRpQijXG5WRJQ/cKT/BaK0h3OV9wauy
ilPsvEMjMTbsdFub3amxBA8o1/jclbYmw/hnIBfaF1HB1vwac+X3eDTrkYiVbb9y
ir86vEMIcAaCNkrwMlSLs9BJ10ojT93uTKNjfLNRbiU9HsqZhJsk02x5hxjw2grZ
JFSvbhhLA4iAEvjz45D365AZbymdthTX3ej0U7hqhL4q1cjSNstc7Lx+1VMeLidj
CXLx4JlxrmaaxJe65ZKFVkcC8/cxs68K63FvJInNu4gOsEV8j4YkGD/KCPpRsPWQ
1VaawYK+nMzjhmzCQKHrADlpgiaA4qCrftK+fl57BXMLC148rM/ZE3AoN+h/b6rz
8Qlvg1PebjuSv7fXhjRrlYTo+t3gtsZsgITXlzcDN0Y1alXN4p7syf2R2CitbOjM
/cFRPzL+kdte4fHIpEWh0DPrjHksDZT1uFsBwS2u2TiC9Ux8jgUo98bULQClE9S5
WlznP7toe2jHWMhKwMK1xwxdif2zRqJ9o6nySLe+QLqEVSWzZItK2PFl/IMmJGao
qj8w4fjg3+YwiuZJxE0rQQ9xF36Owr1P4e4g2COejmFgkODqRK/Xv1aFgV0bcU7E
dhjiUXicPHVUt/Ni75wFY5/2C1u+vKcheiLkpuWO1iZjWkAFVjdh49aXLlIjL8s6
AqhidjNW3+UnyBIGabqTLgGjpFGPEU9aEcNJphCtxKQqCB47zpo/eK6MIpqDoTdW
yxexgJvonEhpg+PaFvhVqJx0ZQNqf40D7d9x7S6YdJRQVOQMcsmNVOZzhy2+rqRf
F9ybuQlUVN+Cj2cTWm/9R72rnAy+iBBLepPZP3WjLO4DpQUO3M04FLdRfpjU9d20
jG6SAKrjonTdgnnMqab+92J42SqKvoTBKYO0C4gLpgcynKmwuOZGyoZ+wF/XGmb/
StEzHOnojHJ/H9zY1Gz9UOrOzlpRS7dDI8HiwIexZgqo2ZHS0nIPC4ddWf0bWdS2
FLA1jxVVjyuGxQ3nUGRRSuKr0IPN4tkv694oRVPa6oTCFUJ3ORhF4unSCOB0e49r
2hY1prOGOXRYhs9SdYmngq4UCDKIG9ZSVxT7TK43vosBWIf0x+r3SlRLRBjYN4WK
xC2lxA3TxoB+JqEMfkKaOb6gnD/ULhB1ETBv1ikrfLkzTRGZuLjyUEBr1zjw9FOr
NunlOnwJCCmMOAaSsj3EsYWC1ttsF4zpDFyAG0ce3k0Ao0x7JQf5jfDl3thEzV6w
rBAIh4mqhueE0mq/LKmedFVEMq5rGOadPDPjmpExbe9VJ69Vr5UtaxI+6HbyzJth
DXYWRqH06BJ2sJEkHCOgRV/nbwYsaLU/wyeUPJdIm0C4jFqoX2G/z0GpY227zHwM
BFPCe8PoAlTDt1QWONKDkBMBQVkYs+gHYaZOVrGqTt0H8dIf1IjYtLFpkpx3EIil
AFNl9DHg6w+mfLoHBM41U0OrGoF9aSIARa0fEmIH5iYl5yTqfuRAGu8HCqu2J3wp
UQAO/U13LJR7Kfa3khkWAhJFAm4vtnTq4K+Awiaa3S1qzHqnu6+DJ/U7Qs8ywxml
NFgRL2Hz989Ty6lr2epLdRy4VlTY23I+oHAlqENZc9B+bwIq6esKe4GtyeSgvL3u
MqURIZmlcmOh2ZpDzQDzRElmGW08AKyVdmw4qIOubmO2igRZfNJWzr4HVGi70iRt
dQvWWr3YgaVMdm+sjARcEBYglgCf/phuGl0BvELEAcXHgGrTVVUQm5UrtOjjSYvO
BmSpm1Kn33r29GLRbZI2gC9rU/Y4MNsWs2t2ol/O8eyArrveLjkiqKxm2YV/nKdf
JkeCcRseQiBJtjyZL3YY8cQQkVpLQV8thh9VjOfwGQ55e+r1xbK8bYA5iUvg6OAp
JKQRwukOt7KTBZRDm8P0TtVZo0Dcedbw+nE4voFxZRE0S7YMNRsvyD1cp0ZaGrp3
WugQktJkPWc3bsOSCq9qpQK+T/73V4XZEgnIajDrRYs=
`pragma protect end_protected
