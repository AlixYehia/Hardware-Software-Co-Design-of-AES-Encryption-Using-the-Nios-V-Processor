`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TOpgwnzasohT8s/aIGtwkEBY8Zi4gwX4s1UDdA6LXpkyiu2YcKL541RuG5/4XeQI
ivXGpb33HgcrWnxt+pAqLV0Hglqf+ON+hyvE16oy6wlLzjGeQv9SPI9PFuQBCAmI
p0mU8KwyddtcjIQBb7xBzSo30scqrlDrxgHhGaQyfmI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14272)
b4xabfQ5VFILBYThOlrQWuxM+hhl9OX8tAHNbv8P6K9wAX/DfzM9m8tsiqi+I1l7
5SuqokD/h0egLd8p0U90dsS7foGYjbfABagjTLmcIZJGU1Ho3GnwIZFM8DrqOhzu
lH5skjdmkk6t0ruVhWJDa/5KKlguIR9TGZpkr7HlFO+OxYMrnVP1Z9NolGa3taVs
SA+lgka0VEr9L6SllyFq7yg1L+tg4DWForack1ZEC74jG9h4H6W6nknWnKCSl0W+
Mqr+ZvXRH1rNwwmmP8lDIhbEhAwxCiPIuVGbevsDmcbD0UZsZ6REtSRfstDzOjyY
tompufvhGHfbYkfZDx6cpJNSHy8WWo1Qmao//4hgZsI2inIx73BeXJn7HivHPdo+
0PWXhKiIOlbQ0PWPYsJ8TNRJecGq1Ijp/flE7QUUiEKjCf8bJsvEbJcOLA6Kq/AK
2j1T8nPPnvx5AEvWmpZ+Z7YBUmPdPzswpaQtIm1kMq01uQnhV/ryTYp9tS7eetul
NK7V4u9OQrcOgx9IDEWZhTXC+XGNFdSf3xQEXYCnhtE4MovhZMLTQe3avdKGBC4b
HDq2Ni01AUnjcmXpAYARiFKq1gW+i/ESfzZKRXkhkrJNi8U3pa3N+QJOFpuEuWZa
JvyAJtJDiIlxMBoDUrgMYHDr3jCiAQXNQDPkQxiGIiDP8PK+TQ043VcMm+zSNkAG
xwxrduFEvkUZ/7XvMYlLHYi4SraEHVn7i1rHsDkeuzU9o8ToxcUWoT2NSe4U3Yhr
Y4qPfjP6+E7LBkWUFakw1wYDIfZi4aW0FjBm7ef59aMCcpEtKpONIb6Jbd+nBC05
6DvYGqrucFF4ZUeVgLdyGiwneP7MuKr/cuu3exMzoEtmcWZxkLXP+UerX6mNgwUt
Y0nnWikXjxBgsXWpNdnetwAU3pgIsB6AMqBXEu0hJs2lMN+QM1zpvSnWMgNbWK5Z
S+DHrGlUQO/Zm+qMBnR2IrKSI1wuWSi1redodFiEzrRaesYc9Jt4p9gJIc9vrSkb
ZA3eN9+rBvIuen745qFF6Kn8yyWdOzfLYyxMdLUrv5YxU54HpyqThp8c5ifSkzSR
ogaugvt+eyc+QMT9dsgMKDs8VEIAK7Vw5YP0uH25OQrs2bsRm8mk1Nr/lu7a5a3R
+hZIQ3MFSH+q0FyvsQ3xRbkJex6gsvIRwDlTR/aZvT+DwRrXnicYXZv6VL/0VQKK
k1xPvrEQ7H25/zllAbCBt4Mr74Hxo+Mm/z6tZ+EjuyaGu9sZMuUBGbPcumcTfCSL
/r1JRIgJlY3Fvx7BLGNWxdMTEfdkDtpKX5TPUjVp+lDivy6wMp0Kw3bthK9mEmUp
pATFD09zy/RnP0AnVyw0UGrDSVuY/ourjlSOeQx3MBtOEOF/IZrFQobrUNcntX5T
MbvCbIaMWkXF2VKUKK/X8Dfu/l25a+pcaQKQPIbjYfJOKbz1VSdRiWmfPWvlCl0Z
qerZ4Z2bMx7UmxYaeBMX5xFvSZ8+Js0yv0SYJqwXfHzv3CchghiM7x+ZtVuyFYCu
2bHWnL5bfmHik2ajdEK/uCjNzmDRp3Gv5WMQjrDzs3hDRdn87XHWgmbCYDnyySfU
277uxoj6TG0x2655Z2GUdtxlbdFpq9Nz/gBmf+NlK/43Rwa8d2PA43HF+LEkEYj0
E0PeoKZUJ0fM4KOw9xBSPKNCgKKOq+oVrIuHCP4EgOcR+ifm8KYBrynHJKN67Te9
quGcq7HZTyztoQKiBhneUDCrrXJ20OtT0VAUvvLPBO55y3FwlXGlMGRVqclTthOC
wh7WtMsrDa6s/puDUjMf9Xj3AITCGRJvI0GtjASvNGp81iIYYZKgRwQY9LwHXYeQ
Y/z2qOV915cXM8bLPlQ3Bzyhv6HJOICY28Kz0xQFnmUH55CtDr4Ne18ff09bsiFM
GOWIL6dSdIq3Ydq63ECUMmaw0BSuoXDSrjd6VVOpUya+q++kkyMZL7C8pAZARfii
3uACydheAS4nw0LDD1nEQUr6Bp1f9VWz3iwM4j/NWtwyXZObrF15srKA28X4T1EH
idffPGPC57SUnUaTb7nC4nc0CtolQvPiuEf1AsophOnLWLlByw4SQYPoleq+gyHq
zrp3lf2CDK6MhpmckZ5xU5vM13xrdRFkizmiPElgkvw1TCCaAyehF+n6YSJFseV8
KU7AngiI+1DPbMmfsrfK1lX3fcXHQ261gBFAEX8rh5CfJuSWB5kAizm3uqfM+9rt
h9eiZjo6+X+uw+k5lhdYes5sBq9A1e2Xe/qdbTz2OdpxTJcBOhHICmtghtujqeZe
jWd2lqkKTvVzpwL8Y8VOXDtz0xUnT8ArA71kFpX8xzCj/n5wgAgMnS+lAkcHd1wr
pwbNSp7Lfcc38WnApc1bWY2aiDsa1/9G9DQ0TPN61whBHzcW4gNHqKxep1tHVgM7
HXDUpsEc0OtPbmIfApcSP5hcn4psjHdrT1dN+NmFv/wE27fD6SBcCkNWabDvKPrL
T7QafwhxXY0ts4H/E5mwSF678xoE1rBAQ8p3/Cl/WPTtpXDCbsu165yyjDIoSqPl
3NCF7NoF7AtlvCZ6g/6mhTlju9eaeTT4fvqOe3RC1mgfeTYLtqLO3dp3SHwTjx2n
Hrqn0+Ylw/dBjB0oj3JUCXO0ttYBsl+zhcKZs97PyRYqD9HRK0t1koTC6Ignpys5
cyIvazqHEAIPe2vA4hvGn7pWdv9B2pYv1tXM6/X2T1ybEdHZzcK+TCHVBK0ok7mH
6t/18ZMBFe3HducwZChJUF0jiPGjw9AHD/qRCCkqIHsUr1PI3cCjWFf/rmnJgEZb
tENYedcJwhxMUb9BcYpx7DGodWGfFZ3IV4SAabkr3s+yfXUHzvvRPP3y/Tay/EKS
uQ8LkdHLGNf4nSIQs+AAskzMYhLdIHWOUuKx/reyIL2Vah8QSWL0HQaLLBDTcBWD
uraJMgegx/tffqqaYNmLztjfXbdneXPO+2NRZx/bT0DezB7FpQIq/PlJ+9GQw78y
o0I5ff6QRecw+zltFLllcMzJtzen3ABH5qWOyJr5LGBbS/M5YoJTP+ecz6N0puJ6
pghNOCsfCcKN45GeF+jF73H1ApGorirjl/4XAlZQvKQO0R6U7++6O+fGB/FZXjqa
htQkpWXxm5cDFE2efTOfKVLF6oNtGWgQkLVSYkLNiOhqNqYzNx8mVxtdiir2w1AI
ZGFD/97D+dDCcb1YRUx4TEsMGioNEP4bR7MdoPCH0Xh/ep25UoavS1AfyBoEElra
FCYjOPlPSRcCLosDV8wjHCQVmMAlsly1pzpAhPCb2rFWFJlK5LcZvC6RbaMCaPEy
LbZfvweJsLhEHE+N4x254wXVP+XDU1K8cfqPDtKDsAbOejbgaqScgS3KBOBZGbUt
pxdRT7atx8+nS7KdZzwLSgtS/3iCrEKyJ6iS0nGL+rXqfoinjZWKdImik/0jkXt+
xE1FsDmNcJj/He3ButEweSsrJnofdv82P4gJhMebiVQ1qM4Rg8jtO6HIZHmM15TK
PS3ZqlSVXDF3f7D3dKYwonNs78n4Imud3DHrKGmhz7c4yWmlXTuWXWlDByK2m3Oz
OvNW/x5ivBqfxub0QzH36Sm71+lsz01VbMxgCE6J3DgPnxCQ7A9dqWX3jo791Tg7
nLGfddOUARwN52ZNDYhkoONy1fRsAB8TOY3CbjwEWRy3LF9LP+tyqIJZVC0f7x5e
M9OwSt3t6tHl042shQvH4xOwgMH6vaEMeuoJ/jG3ByJunil/iAMMNKJ+jNPOFQI6
trpH4ku1eVpaCUvmP1UqFjje884WSadaWtpVxTS9G0WfJVAZ6EtVNcxAU0AXVXh8
wxbwEgftnPIdqTLev4cm5JRLJqCXud7n8cY/1/y9PTK3jWv3mszWHIrJinE+hO3n
84dSWENVO7DIwMSpy1YDpuUHOW8iOA07c/1ZeAMh7CxpJQaOkVchmlV9PbGTjnvW
YhywBZF8/p3jKu4jvMXjY5lYMxKjgEs1festxw0FgnmTfUPE+So+HTfWIHt7zu7O
2KS2Fn+CYw0qHlwdoInkElQ4VJSnzpde4sh/BDXe6H/qEps0PzI1aGj293zNAZYB
4afnL2eX263xbTM1A/eeO7V6hPZuotLzqOwHLfyWPCy0KIn0UpwGPJmrY2crlicy
RF4jj/8BVtxO+XHOYk9vQhHuZdFjOHINPj2YTNY/HS3FkrYCuQuUarGP4fk5I5Yg
R1Z24Jaw8XKmzAk5ZRhdqk6mkPXlq5RjxU83iJZSIhfFUVQ8niZaJuCowM3oilXs
XrxqBfBOWZCNJKVOiplViuYOjTpwkmpdIBe9MJ/O3+FJQ3xmJEoUStbgvjKgThiR
q2InwXcg9TuU69iu+OV1uH565zNuHXdyCv8dGqAlgsXzYYrgAkXmlCv5PLorRbLT
dsraPmsqKC5/lcZ+YOc/fQHdZr7kMjzVxSO2CYj+Z1I1QV/tup4t7hQRKslNzSIg
DFrbouHZLiFm8084JKhMc6JwWitbo1plimV+M2+9xS5PvJYLmIk2UbfzBwmc0THs
1Uzv4ymBn6rs7uQqiLStvNrTtLnkgU3x0e0Z/VUKgoCUcRS1XTf0Btgll0m7DUQ4
bJz/LH97OSIag9Z7UJjUaa9e7RieUTd9djiL6GtHYjrvG7VcoVyqEnMB+01eln4a
aF9j65mNeusvMRsFtFBFpM0MWInF4PNcCPF1ILjSg2DtDYc+PfpBK6+qxvDWvJXT
gg4X55NYANfF65hrIt9/ExmXNtKuCbX1KLzCyvLrCo4qrd8S0F+E3dYrNKdcukcc
XPwN6m98nuewSWRJRIhvUbqaMS3YyOx2i9ohDzEisxsf+aW9g83etaEtFusXnlt5
O41F8zFmVBxxu7THusSraZZi93kf1hfcCpncyWuH/EY8ba9QnS50cqFm1qOj6oEW
Fkyn8cXRAPygHJBpVgX5ZoNRmh9dDbRVUpAfAuLsmNweFu5zYIgDXIer2pJzPmOs
KOyCR/qekCfCew8hu7F41OAvUM5/R/KHlZ7wJhNKiXYGzH7NQbIReKrpGhPiMRWM
YrtFbHrtm5BFiuq7Gv+lViZqriwpU2u6iziDH7NG0JVZMNseaYUcI7MFhyfaqabG
L+ss0/qd/M0iGT+gFbcBWXYfyeHPODVk1CCW4XagoloX+HJlgIjkym10hQmpj5Lj
Ekzu66VuWpBDOwrZTtOQxfduwQT9SS/Mh+2AlC2P9cr+VJR0lEgLHgpR5XjiSkRM
QlKVZKYtVn04Oo6ZCMAx+iVFlp8NeosVDJ5f09jbWp+pXRLS5vs5XyLeqpqChOVd
8XsIege7GNBhFphiFGcojctpkSVKA9ldbRNBh2nuAZoT02hvpFO5z7gQUwgZYucf
n7BwVN3YaDV0M1rlvamTh+STNqdInQ5mJ8hIlsnQeJ7BR7DpQzbUez/B4SADwfNW
l1JavZ0A9h31sR4yg8e9O2/SOLKf0eHBmEghkqgQvjb3W++rMJD/GnYbdIPp/6cF
moNVQWjDp1w5j39WHImbwnt8BhwD05elgGjxszvvqkMebsq63t+rMQwCGAKLhX40
TLw2QCd3c7Px77aPfV3RWEBav4robXY60S/VptfIdLcfgzhFnvquqfBJydFB6NQ5
AsmXlNhMKHLNIrJH0Qhf8UZk4Whw6tCX1CJNchRra3AGbPuz5VXP//SKvorRsUUt
697u6f/+ALBH6YDSD+YwUOZO9xSMKkc1jtbhEvoD/9OhJ044Fk8fbWrlxtWkvkm5
5d/iwpMph38qyg9HhMPKnBZB/XS26XXizxuEUvtm8Q3t+bs6/P6RhrPIfT0dtwcW
wIHjDp2j3Uz/bAHsUKllDjlOrU02pEfZFRXEXIoD0pUqZWw7lAbC4DS1y5iqkpxI
/PDZcXGN5bi8KMBZm2RQrZE84RvZhnCPE2jKnDjm4qOvwZS6WEne/OVnsTpnGlY8
xd1k1k9LiAQB2B/CpSWUJteRNjGG9s9P1zH/EQ7RrNawROM6IPweNyXtkI8gmQBt
EBxMIoFweF+lg5ERu4uG+/XX6BHOGtwoEvqVMopcfqHa15OLuLl0QIM58x6Xw9tF
U0whapxqH5O/a3LCwvnztAVC4ekiMWjwyZDqgIfzx1SqoePqdJMI3t0/LK1cHewV
ICQw9dFjD72XJfr6Wlg6nmkM8qXS4EkBpbjf2RgIygHqMEJFwlTV7P3LkthWUvj/
U3439Wc8iU7rkjlr40JpaQiPuWYaq2szy7E4UEBXOCwbbMvg9Esu6iuyFcGLnH4X
/mWmjZKTB3KBFkPLYHho9aKRXN8Roz+isNm6DHbBvViYcvTBIBCtgftaaMq1xGsz
/lInKS2v/F3/xoLZNZC8o9Ys2YoiiY1mYUlS7ZIBifAlsXm/tEih2w2HMEnDSRGD
J/nxdDX5ub1yBzCB/VAeuoVaHw6LzC4M2O/eWsELmF8gir4ihzziGAj183S869Z2
u78obMrPRz1LY2iHThuBQav7qzJhvCuWjTzuZ9n1rOxbkhMY3gjUF7Rs3EaDKrg1
VDNOxEr+Ny2ww5O34r7iTuAHpk+508s2HKtk5FhBjn1x1NIQ3cVWJfPCSnV+BYok
WBhaNqQCUHoDDa/I1b/OFJt3VIHfIl9+LLwq5KLUEBlmHA7QFgCV1HIMSnSsI6Yh
A8xoQmFDOfUnilzVEL1d7S4+Jsqnw+h6EpZ+90TqBg/x9ym7ifxVI67767jJnVWY
gcWW/9xplRZ9JjNfkc05loIZ2iNC8ng5fCx4gHcfKsC8njoJVjHG9FkrMG7zPcQJ
ShvQgjGv4G6LiDgGGuLfxhYE/gnulxkO/oG62PR0lysj5eM4XSwWtOvjqwh6soqa
G3ItnDmcjT3M62DwYgXMw5MeH6d1Y7OeJKXMWwdD0ebKTvQ31P6o8KFpccdSjMxz
+Pv79JAduDMrzo1xfbrRJqyiJuPu7u2pcPd1Xr08Zv8gQQdvrvaCKLKuE9ENEzmE
E+hEnyJA+jPguy1bfpl1uwJ5sCV/v4bhjZzp5Zw/d0B4PKsr6wHhQbnv8D4qpLkL
iUiRZjrVEHhedgXSl8EbjhD01Hws4CEQr4wtfiFZueyzb42nlxV0TDleo0t0/Dmo
c79bOCNUM8dbYiFzRJRAcJk/GtSc4A8+O1lhXeEop5XPmYOzYfvtwrzIPWmUsA+y
cyf5xsi3dohBFgX00/KvZTeJd754bqEjuNAfkds9UUfNljeVklnTU44y8/XniQHx
eym6+Yx5CsX2dsBA7tipTMwpiOPaYKjK6x3BoUh2qKVFVjxpL0uqOSrhb7XZZMO/
FIwAtTNsG+R42z7jqjZYPl8kUNyVXG+CIer7sxYluzlIzG3cqWEuDgTrCFQAAAmA
78/sHZuAw3K/s68Pw/HDvIID1QHpSd64QmvSsb22j9m/hwXQEoYjLOtCGxKUe6Kq
6tSaRUCJyWrl3DBdZmWlPlIGe+3OF+rhfyqRQJejtC48S6XjNgeGE0kf0BtXatEl
LzSyM0JcsLDfkAV1bTNsrh0EznzzSilUJrpScOTZ37LpI6Wodis/BsIQ4d2BLlvi
jBfecG6pPWO5pirFsu3mPjPtM7TrP0Y8SorF9ZYJLxdm8vc0y+0SNgjCUWaYMLP0
h3Tewfwd5rj4hOI7dv0y9LoT+B3Nb4HYf/ESQAkwP4htuboDeuAnJgPlniS2mms3
aQOoc04B/bhTAAsciAsPYqijGsfGW/BoErDxoiE0tVmxU2/bffQcd2IZDpMQ5oV2
P/qw03yQVbq5bWAZoDmzUTwUFeI6IZRPrTGYaVn+8uqDbE0reVbTKsCvWr2/ZKlf
Ok75QxuTjlqT0jmWl2orrD84KVJyQe8nLN+jGy11xtGTvp7VdMf3CPM/AR1BZx+G
r+bwDDRnfgFiAEHYFMb6wVQXe9+UnKCD46M8bkgH+1kajh7zfQXe/fIx+9Ofn+wX
bRkuOneuhw41XO2bhhK7BRShg76yDhH25LQXJ81UbOQQf6moOG7kmXSpuPXeJywH
sjN1u9opUn2H08sbH5hBXjyGXg4WwfAVDtCkn/CWOGLEsgRhZd8h5EHbqpUKpxuj
JMHswx6Va1wTKW2mI7VHhkAFuDbReLVKQgUrZEx6xUzOGypoeemdcRe6+H5H6jW1
s722s5cWNGGZjXrcZY85We14bodUjJQlMSx2lHZPVSb5mBo3SUgLHBgnoOr0EIQ6
wPHEtYWaJBHGDf2WN8dq0tAPGTBDUI6a/0iKubPskRochNafgFKLNtb/Bc9+JHPE
SNapS6NhM2eTCnr8KqosRViUdOXlWL2I2dj5YeB5g/JmQi1xxTOsqL1+Mj92K+C8
MGqhESM8P2uQ1rauvCYeSo/bhS0opDscIDguVL4g27YP7501ugDVf+Og2l9sy5Jh
+0wEZ76TbF6jxqRPx1H1AocA5DFqSB5SNoeXrBHxixYhyJhW23yQ/Zlddy+lYIBT
+uBM5cqUY2o4t9y+UqBU6ta4JTJyvpJlFquql4LtH+LgdsWZDi+GMQHBFsK0sTGo
TJVuxtL2h8dhQ4eFJs1fXQEsnpiFqOAmmUNxLtYzg4vBJFcA2aDboGBWufTjV677
CUPrbOkw+H5AzOx+pnndnurUu0drV0CX0s/nQaaQcBiAbg2+OIi4nFk2Sbv8zBdK
jmCwkBQ6DRJJ5dLF5jxFqGqehE1sC9xFqStyEp+8H8j0eFYERfkt/n5LKiDUGuwI
/LwiB2bdVtfu6vT3PmL3faky69CBYdcLHmrtda+JXnZith+SU2PKAvur79Jeyuvn
RHO26fIHliuCeyQTtUd8WltpBa+yOeSVVFDrn2FIM2MzlzgmCV3O/Mw4PjC6/mWW
INMkY7ikr/CN8TcRyCPGOPmfypp/YMY9EkgNbdrgUeI9e+fx6TgczpNEwm4psJ81
L2rzjjWgmhd4p4n0m0LxnE3Oe8aWQVDo/E1f4UYvVldUNRR4JaDkA7VpCz6fUGJx
9xHbrShPCWinFgHPZry/aQXP+dyzvjBnCKbOPnb8+YKrxaKu91mqspL6ym9eaaWL
LNII9uYVIwXIkvcmf+l5tCFrIYDxghpEGQcNPSaJwalCTZNycVHYLdYTmzC2U2GF
Vpb0ct+WCC7Ur/xkqQWR+Sc2NAys5zWgyvQsKSt1HwJtaCUX2iVBKyyImeCvTwCA
f8VyE8T+Hy852LlpYccipKW2lO8kSn5skjLn1Uz2HlOoNUZzhhyFMMQ+FZUFnMIJ
XSy3WMGGrubidQZFjx9ZV3b98HIYr8yAfVzjr4rY9aFEF5/42K/MCjM133tFZ372
tiZVp7teE8NTBIwb2jFz919qIhOHjpLobZbaWl8f/gymv+FGLN9sWXNgkkqYCT59
kDKFCbEDmEf+/IGxO5FBocePqVNURi6RDsTOP4esTVB7ucA/LPabm8rTZItXDyzZ
zTAtCg7QwaPpiqL8WpVDM6wj/6l+192NZFfIrWc1HxjRTCWc2ODpBD3T7esYj2+A
Y1GKCCeH3NzxZTWYz/zMsEID3F3IKLvMUSDW0Ca57xk49uWEMkGzsQP5PHsP8n1A
XSg+X6TFMGxnjS7iicQKHcUKcqXlAdOKX0Tk9dmcZbinTy02yscKe3nUFEk2OTbb
Zus2rLGxYxDLdY7Ph0pEzUunDqIcO1J8jA6J3Q6tb4Ef5ixHuJA65D619+scTWpX
p+S9Slb3tZV1Jbft5V1GrYJLy+hdlWnm8Wvfte9sz6kMhXe4Sp1Vghpo+ORnQeSM
3tNoXmbLXb7Kpg0TVcgnpDj39xrPxdusXUPK7vckqNRgOtz2XJaudtLmsy03nYK8
kp1a+6F2eoZoKOoKDwwXVkHyntw3JE1R4IbHRr5SeJNaOsu4KqO/piKB6Mp8/kcK
rRkaXAd6efJSvkc3XQmT5iTcJ54rBExEpTIEN8cAx98YYw5mCBEfT/Qnp7aP4GnM
zZldlJriW+m9aT9z688mPHWzT4u16lvhuxCxQ4+HnZNiFWyoBVLXlD8AQXnZer4o
ECDzJIzkOxa1GhgymWLboEdoD3UXaOvVzkkPS0eniPrGZUtO+4SrkX09rQxNtkdU
Ws9twR81Hy2Ze9YrzxS2SrpUTZFAi4+8Evvoyr80zO07Jh8uwMaOFnk+NkFxeKfi
vHqxFKdgXvDeP+BAImeLIA6AxrpYwkCuDq7RlrdPB9c0U3cA7NaCpD0PiwTadeT9
VyqoltvAB+xRNDi6jK7wlyFQJHrDJD45MK0TGLo+W/uxzG6ELBKsD9ZaPOX81f/S
vrDz7Fcx3I3jEVKq4B0qsSkY6IwEEK9NjgnJsXICQyL+l8MMAZGQSQ7KGm16bnL1
KNrl7uOp8kmAlFKwoij8jyyrEBYJ60bUeIkFUx9dQrH+iujA7c7VNlDiCkZweOsN
aAfCOF4Rox8cPY5DbHP44CY4GR2/Va0t/10pzqDRaedxUSS5JLkZY/LMoMQm23Mc
7R6Yjp7wWaci6kfNG5ZAn6DeACQzB5HzC2q381br4UqTvA1jC7JCKaUkU2tjE3Bp
kr9ifc7alZBvSDC/lgtTZidQ+r3miXIFBO1emoGYCI2cLZTLuiUvS2U/BxurIU4D
CmBrJrzL+URB6BwDiV80dYHlioDsiEGY18NfmAQ6lwzSpIp7u2ReY2q5cNtPFj1n
QnwR494dAUNAPd5jyXWFDDD5q1j2se2iyKwfphz0631joZgI4o2wJ+SeD7mTO0Dg
eqW34vkCAx4XtQpzw0YkD4+8pFxj/xOj7w+6daf2tygP/mzkmQ1S5GKpWO5tyx4c
4VYkoOPJiSnsWk6QH/ibQjpJaQO6ls7J47F5iKrHLxesxqLjx/IyQSJTWxud3oGo
+8I+WIuljP9K/ZU4lbURhWOfO/Mk2Z5AiaZzeMifg7D1Qr/QpvQnBxFuW5eHkKQv
6bKdzT9ererkEVsQFTox3ek3o4uWitMYuiNMrDLMP7McpX+wb86JdNKnQXA2JH+y
dc+cIomgF9n+18YbI2K31BYgv0Mr0Ww1z/sg57CTRyG77f1y3yNzpVo5VuYc8/FA
+U+9uDSdcaYG5g/O7TdcoB1JMBxpBhYpsiWMhD0/hONr2bfZnUam7sSoV/vp4OA7
DzVie3oMtt00NJJl9DaBoLWfbPOsY9Y1DiMHnZ6fy1O6jr7Q73NDGviPx15gZ/yA
BkukanHGAXB8KVr0E25B3vrR00ASxjYOpCZrFjz+wnJM/tzO3x07AfI7Qx1Uv0Au
XEko3otuepug+Sx71RmEzScNtrevNk9Eed5lnlH/o5Ci4ta2Y1ItqKDCE3Puxzrk
TArkU7MBbw5pxFDCuc2YJNXV9dsjgFF0YU31EoRAJbVVWtjy3DOgstZyAr3C5uwA
vRBHcXYnxVZRbghtFIWVW/mda+HB0MOzmsAHkl/j+oKPlUir9h8DGtoTvPHkJ7It
kOplbVphNgpr0DJ/ahX03mxLVJrHElXuhQe5+9qlI3vhbmZ+uCCXoVU7IoKNpr6q
3DswuSUllPcbJ96g9nFoyZJbnpyoU4hcLZneT0Vz7i2oEBnnKMdgOUwt5n2yAJ2x
aH3GuUrBmP6hUGsXlPA9omYuEDjE15QKTeQeQStk22loAYG+ZEzW6+Jo5qr97rmy
WoIweqxieDVCIKKvTmfTLVMLZgtMtxpecXysIh0TIcwBV5+9x0jSWmlGBZl2z/kQ
52OQPvJ3j3gAFS9u65/q++zRMK8QPPRgBi80+Fg33HFMJXk4Nz1T1/VzZumRjPk2
D1eY4FuLBQrEH2ZL79rEu7f23bRXXkRcnKqBRKd1arq/FUzK/sGCVk/DViQuLQM4
L3tucYfQ4M9jHvqhaXzehbNGB7U9kOCawRed4nnpib50SchDi9ktZUbRj0BPwVqR
0zw9zQHpRUAaql8+0hGYcb0fus/bB6MIop9hLje92B/MY3rlnlQm+S3j00+ib3pV
pstrsgVqabiTEEtej8mtQzDAf7ZxaJCPOPmr52E900Otc27STsV71386/OROxJRm
T/oEs80XZff6UCI349z229tYQO/thXgsRUkFIaAUN+965rOJR+zlVw1NXOlEGPMs
hg9JJDQx65xuLMiI9qjSoydqN/dOriZWfwun1yIT+LLksDieWF6yzofscbxzfq+T
bGGcVPsm+yxY5a7D2NelwpTE1XdHg8kUhx/V6QNfG1p02HEdngTCNeKSsDH2spFA
ZfH94KNJ+2thpf5MF3ewD6mlvmG6LALDPG8j3gHyXeMpKK8U2wBa43ygufDrUvc4
yQJnvL4AiDB7rQaDnG73a3UizEVKtjz8CMwyN4OTUrldrC9v6F1IDOQmBiODNTzh
0SqZ7dOZPne8/VMXE5ivfB4fxSP8XkcOoYnljzGW0c7CfV00KxOvdEnXx54uuNTo
ziBS3z+SWvhm6CN5z0b3g/42qt3m2NdbgtQwYoWhWpsQY+U/kBDrtEnGzgd4KD5Q
OPIzI6GI+E0eF8r7HNbp1WnptR0r+6ZM9J6dlxWxhmBlQqX1HsN4G8qkUckPlTVQ
RX042MwQ38O5zvsvYhuvbERi9GxF8n9fGFQtB2KlDbycVu8qbf3hA5PcjFl5p8Dx
zYVdYkCgtJ36SZecqnHdXBwbZ+eU9xDfT3+mxdv+2bLiRcMhxi8THsdbnTOLc2um
mzF1CF9UrfKAjieKTjRa/dtgvYJMpdUG5UfT0JRixEQRfZd9QjdcvcgQFay9PPWs
3X+vV3sZ3ZEFcBZEf6oQDYFsapiN/3TYooPFhZGMwvZgtxXCXyPr+hpStetYsE5i
dAlSItx9K2FnOKSOcGwRjLBo5rv0ayw7zqphP7txZONLzY12K/Sr+tA/EoJHJmsj
VzvJ4+ldCDay2V6n2XE+63rHual+myeQsheGx/Xac7quozyY81cryCCYHLXzZxxp
PEs/529nxg1hvgkWZ4VCju0WFWIXKxNddNBdlAtcWVrhFWzWTK1cLA59g8PY7NA3
ckg2gKN8bp1AHk6oqn/59lAN5Xzz01erMVkujmjFUxGOm0y6T59jyxfrlluM0M9o
cVifhl0yMMQA+xpTSEfREEj7rT36KMLxLlWLuUbqwmQCOOITF5In6pIjPdR+OLEN
YY6+BquL3MSyIaEE1eo6HRc2vFdMM3mnG4ZmpI94QcN8fkkfgCHhVBXAWJIQhzxR
+zSQ7YeIqKA5qXd1bkR7v0WiZPTgvdfY7CN8bdi5FUctcmI1/i2U8o9W3AVn4602
gkxntcwJXNd6sSObMmzMEHW73Ok66b+SafQpkfVSUgpARpezOTLRUSsVm+qaziNU
KI1cAIsTWZLWsxuuofOcJaruIHmHaMp/ZnuNSaCmnWoLKqXzq2phuxNUGDimsbE5
4YfRxhIKecIpJHLSMPxZO/BZgQVWL4qf7N6xIvMcr9ovUfD8pUq+nWYrYZ+dYqno
kHSiAFCVX6w2mwiYrJrr7BKrBN2zClvzfQcRvmT0aYr7XIkAokswJI3te2+GfUXq
cobP8JizP4JHxrttoe1r86ZQiBw3mqqiawZcc+jcFhnfmnuAwhxlnloRXmngp4Z9
kPUiXuwufLh8g3KgnNI32wXABLH5VI26K0HkWAcvU0d8vwJ+3o6yyctH4/L0P2O7
23hsG7cFQXdajVMGI2zoQBVytSx+EMKGKQmhXwnuuyzYMSAq9vXj0Nkt4/HX41zI
yhI/mHE+Rmpddd+JNO+suOReQ/exoYl/z9f/LEC/rTgfti7/AlovStFgmkV6qNfv
7NVXP9sHctM5FPlQaCjjt3aWj1r76CBZ6nHCcRKnuzG9GulFAyClVzUvn4jhPgvM
I17ztP3x+C3aYYeGFBoalmDaVyPHLldgmvdxFmoCgO8ob/GfW8D7KghZ39C5laE4
D4yZMnzsUKCTomfs4yJxX+S5LwoYGLrj3WQ2RS6JwJYnsTP0TVX1NZzHDF6zSK98
I98btIwuZnsdm82fBKhs+a28t1CsGQo0xr/494JJMySdiFS1uy15VdkdP+sxDgxR
YbnQfMO9I9CLeGq9MW7YlA3SW1LiAikx+LteADXK+yzCSjxRa+TfuIdVe3sqCZef
+vcSSlxOMrwmAmaWLiZeFa7BeZk8MaXOp5VD2sm3438X6S+iWJHo3tJfaCUiW9fw
95jA6smi0PNaVvXzuzqwZPn4eGZ84ejHyhJii2PIp90Uz1Usuh7sRJAPJyG3pDbt
jGz4xlAHXXggtBJjp6LV2E72IrjzU2XTvrF202vcVpwXihWxWra21DjQDWwrqrLU
TqPu6EV67b5V7r1aiHkUUUbpbUDbV0/VLgHy85EDeBZD2YfcdOLa7EJIdbJGKApR
GMcJzop6mhGMJd/Fz676UImckizSuaPihYk2uDLB886tLCuNbIdZDPQ5z0eDg9Ho
Rt4hDhWdLFmYTzIcg0Tj78bqm0kU/S8ylXjOC1pGhZHpc/zO0PXRKq+/BTsY5ail
rJrF3d6XcyTuUib6BsO9ym2ETlIHKPD2DcwnyALP5xotPX4TOIqngI1w0RE8D61m
9DtP1Lf2Rc5V4TX4UMb4dSf/qRCrMJO6iKFp7rwYUtQF/5RaY1mAf5o03W2Tyhv3
R3mRzbbzkxlD+IFAmoGZGWT3ZP+GzbRTA245wtsX8j/Dr+a847A4H2T+XA8Oguek
/hl4+lYdkhuDp4ogBhx8UruBkSlCzCHJMQCUt9T5JRCJG00dCge371mjPLngXD5n
FugFQGkdWY9xQuWF/1+HCfjLAMYonDo3dmhSiedCNxiRffL5uU2il7G1BOe2eoRt
11fU7JHWfTQiyCdBVuMohDxE2+sGtOAcLMld9eKP6sz29H9EAcZFbKeld5+F1xZm
MZ4Fz8o7FhGGztbRrXw1Hf38zhS6WmZV75VyHMDuqI6p/3YxM0x+Yg1VD3LBtVMi
tgM8qaisujZUIvTR9Xp+d0tJXRp+CbklYwl7H3Zpn1c+o2hBm/mEWuFW64EiBGeo
znefYcmXF/evfcBSxwM3KvaNka/guWEF0ml6PUqMNsJ7y2XgL8FJLEIL7mcMVE1b
vIQPedXeO0kDMbFsX66iSc1dqG4kzCz9HE1rSdHCAlj6EQxUMVab0uvS7aWk0bpl
PVRskwda5NkvqqDKmhGvqgPd0yzEMnS6WRLv01vl3njxrfOGd87TJbY88TDvZ1yh
ZmHSLC+BMqaxsxp1R3fQig7cWAcnwucbfdjzJPKbLklt9L3N4nylbcUh2cqzHQTe
vk/AymHMJyP6uEZUwIKfEgTN6xvFRuPlILpwb5/8n4PwAJ85gL/Ny2UISmEnNc5S
MdiPQbFHMfkuvQmzTWW4ssYNVHgwrRdIlVsTQ2+w7OL1I7fN+8tsTGlvMVf6Fks0
JUOaQrcSuahMus/OxXi/NtvVlHHudBEHUkIKFngAHQ8htiZ9WL/l2lG5xyY7KBDO
NLx8H33IBXXKRBAaXn0toFLCKozUFwCdG/q1d2zStI3S1llyap0Le8Y98Dm86Ldb
eZUdQtqO2sq5YfCLRFIaaQHTsiKhGUfxKp72A/oi75sdjjZtV3cvuOvXnFHeo7AE
cIqKntfQicMJW9cLXHNkdoBxu6hwqndRaqittOmSuNjwBgPDojlYdfvk8IGZT8yh
x8GIDoidstOYEfpt0oZpB+TwodTDJHEI7lD8XEl2P1pxx7p2vSM9qe++ZTKGS3K+
kNLt/RTbAMOqLKVZXgJgDxlXoQi9zgI068h9FJ3FHoK0+h/pbHXtDxHo2kPf4F6K
yA6ae18OGqtTtAOMjAoUjcs+4LeffZ369EKMY4frNRu/VhtNi0yFpkHNZnWuOjFu
uv9bA21vaMtl1iM8K2cklh0OsGtJq0Wiw8GtavBuVLIoeWXpyJ9y1dEJJUGxi7zc
gjLjKfoZyl+k8XxzWKFvT3n4X0QkGyfTWoadau6CpAewocWm8wVDieT3HygC5c+N
gfZ7NEnhgmxjpGoRYIeZFL7UZTr5Qi/zy83vlGLfqyCQDPKl1S+swrvr9bg16QLp
PkVsasZTjesu5D2ZfxVnFD7o21VdFazu5FCUn5FF1mNzMtwhLfZCjHKcYOZG/7vH
X2IPaqVXUvwlxh6JvDSGMNXEAQ3kOjQ43gYE/W0KNQ8R0fzbx/RW0rA0cPBQa4mp
wWppGdOq3j0Hiaj36YVHQ9z8/37vjd1mY7TLq9BZKr/Yzm8hDcblYhGm5ISe/ntj
44aMvA/f7502OfXDbO9V7prpndcaahO+AtkqXPqY8n+vkdwzv8KGqieiVh9rQN8I
yzTLRX+Pl77Hfbv/DF+i3THOVkLtC9B1tInXaoQB3aJik+aYY8NCdRbnLjtzXiV2
FPYnVKP2+nO6+hAv9IxJx5PCgMi3sct4ahydAI42fFmzPZ34qO9WKwZ2/RNJfZO2
pSamsEVCWrYMxNY3V111Pzk/dQi23cTd+1C4zThCMhpiFuvyuAHqCqZQA0D/Hy5f
XNPpAFIXIrAe4dVJhdP/cnxdCvadBMH6z2a7yjv0cYdMRKxpIPtLqeEd7Pk4DWv8
DxQAD2tkDAvmjU8t9aVjqQawzHTVYhLeoW0tVpyU2aHiYRPkdkGdJ3lsfVYFocC2
AUIRRWkU7AeYWdBivUoplvcyfglLyRB/tPaq0+ppHS+cA88cIM8CFFoRqC1ppOkg
r66rHD9+8Pnu0r55FH0gn1la2PKOe9PuUVXn6DjudOz+Y1yjFMO9mZCeo4iaqMHU
y9nvyPPI0R94eaM++XvnSk/9g3WDd48MBUPutXSYc1Z44ujFdZ29fRIi4fb6+alQ
8+dsCxu4qygq0BtEyIFk1grxMIGQGTfNj1E+ojraKKjB3G8rClfbZrhqae+UVp5/
gSb04jK2gdCeg8HEFgjYm4OGxxOgYXXCCgaEqo9fDbV7nrkH2aPI4VkxL1tQn2Pp
C57tx8AEIU0HcNSx0HknF4eYZ08xHLk8XxJmaHFHlSfVGbdETZ7GWcz/Ik2uGUdh
v/QqGCFds379uvMCxyZLf4g1C+9vwTjrTT6Xmpc0wuMrCGAQsEbfHhCgNh/AlgrM
q8JOSKFmWxjz8wbfS14YCA+aKoo9GxOCN1ssaopyQAo9g79JNlTRe8wvnJc3eJgn
doOvYChtAMI8h5WDFZMNEQwOCEj9yRZFnpfTH3GKxdbygVEju0vT1L4A6VkpnsBr
X8NELVA1SqQ8jqeX60F5ihkGf0BrEhnAsCQ+V2U/YLuoVxRHDIi63F/yZNERBwgw
5WNjjD0GvXN++y8e9I+0OpMQO4vbGbTNEKmJLBiyNQDmtp2OLqlV36ftLeco0lV6
7wdjxBJF3gfwC5ctF7Pk66qVsFEDXF+q0BJ2SVwsIRG1QABgmAwEAbS8JjGmxmIh
Rkl14GZ0UpMZLXCDEzCSdWZfoIIEc3DYBgnXsoEd/CK70zwsrj+y5/+6lj/HgVnd
xdwsOcDpPUX1dFQy3oLE1VZywQOY5FJvrruinMLl++GKOcywQykm/mtzE+U88ixq
9ATp2psemG0DljBKFNnoZvNSgaj39hNQ7sT2fPN8jdMOJq5bBZKYyi2DmRXaAAOR
6OXnKt2Dz/JM636ZyHiNJPWWwI09dBo2KWq9kcMTHI7DpRwKnxMzx1yTRhD+pSyw
DPk3wX2Z0eQ3yOkeQaN7Rdd+r6dQKlsCCmeMoqtdfO/zWQR6qI5QFpm9q16khTXU
dAOIktYRL0RPSYrnX6TjIy9G4Cx5aTjNhPZg5xpqVHjmuEleXOF99fvlOJAesKGL
nd6+Qg/sfPOcOIwNV8S4FbpGP3lz4jjXRFN8Fzsf/BW5NbVMJWYilIxlGdRW3waA
PF/Jj4Ui9CQeaX+joKUmGoifwORvCUi9CJSAxBDzUw7/g6F8FBUeq7YVvJfKw43l
LOoQLf36hgYUGwuL/1rl4r6haJfyXlf8D34GOZWUclRAEBIPTyb02/x5BKdfgpZK
xq/92/30o2NMSCol/5UeVTYl298vuWmTpwBZNCRvWf6ONChQaz9lyWg8IKZE76re
UHmr7q1it5dcmTKV4LcIQQ+NTvvKXr3yQ6UtytYtiKkpgRUtJ6wZhtB3ZNtqFcXY
rj3dgzvmz2RZ4fwWa/lRRGLIkY70utckG6boCV3Z7MD/FSx+cO1RkI2SlmnKW/Vi
9CmfT4IC4m6O5iVTiaQK5/nsSSdFCp32efz35rrb4ZQxR+G8iEo4mNSGjMUAZmlS
wpdWYG+RxXduUPsHktTAEA+srIkXdiGORNRi+SNbJC8RenCbBSuKvSpt/8LZNLVc
iQHWN78URbPJYomYtQt+Qm8LE6F3rc6XQhaCyt9XihjXK1ywqJ5E3hvGRKPDsZHk
UrHxZPNlHKYEAv8/smNrlvoUopfK/AiZPZcgsZm9gMYP9RkFF+5BkQPvjmeSNQJ8
v287QFsB8mNK/7gG30QHEMkEbIz/LpUWHXeRskEUk/2ngDQbEpRU8YDkgRSLV88s
Cak6+s3Ro0qeCdOVRIBmr0RhL4UlMRcoxP0gZfGB3VEKQtjkfrfmeFPQ+aHCFjgQ
3JOxDv6K/BSTB6AkljivBM03IsgR4nO8NMcwAEH1ywve320SfzKpqAOKVJyiCbut
IjHcIuFA2RfzYNNbAvBN/fhxLU8Jz5nFRVpRmNu/lQREkZ2lavx+QZWA75lHtf20
GJJ3EknehQYE6XzFw2CyBRFxTLFOmNsyYtKrIAeCUsL5d8R5AKh+glurU2plt6py
H4vzhTpPfVNVvIWxkhc4DFu0vEEFx2tKMxxzj2k2I2zE8h57aLmDtX7ZzO6sdZOw
FBFkpbnfmAM4hclogfSmZsz2sNH0L9iFqVBVNsQNq36idj0zWQDzjyVrOwRZhP8y
uxfXKwyQilxB34+ddp9eoaCbdFlhnHqA0ZIbWKHFE0C16K/0Bh/XNixLXA6+o9CJ
YdukLnUQzPTe+pREi2WjohkrB82PEKx6deneJDOqP8FGKv97f5zZTzqrD9wmjcJk
UJbIhzCy0Tg48S8pA5qZUvJ9/Ua46gsGNKONz67XEUbwn0FdONAut/0pKwLwhZUq
hxWOKiz1Z8V4co4cOSnsqbYDQ5FSMob30P5eipGbktx9zjckCkPFdcOhJWGRn7WX
pIjWLRBltdf14ZUccLD2Sg==
`pragma protect end_protected
