`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EM5gSMoOrkDPto5MASZ5VYjKftTJG+0HfldHubU9CA62N2bwWTrsg4FldbY4kUVS
iU8exKVAyU+zmxXcSbSuN0s1a4PEQRDRl9aOy8MczNN5F9pq3+M2jJzfVHJRAAWs
jacFQCJTQiGRHQm20EEF6w8RTTITVRtUcXRtTZ3pIGA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3856)
IKKS9sPT6nUmvzoRt/X/V8blZmbFbIiCI6BAKALZ3CgWLbXOk+pPfPryEzD/zKTn
vxy+rFIhuHEO7byJ8CZCAiCQli/R1J/oUgY8rdSrPmoQOMO3QFEOaTgLIEDwqKL4
0HsZle1pMAq6eCPPGxS/M3ZlHq/2T97egtotUe8syXXh93VwP6suxaKAKit6GgjC
HiPNwMA/s/OpG2WX/4Ojp+KDt3OcP+Z9eJS4vhMML7wpZMHhjJdAAeBucSoAS7dD
7y139brmmRJrG4B8v45ToOXeit2oyQQrr0proClNDp6TQCPGij1PH/g7c9llp2ne
M6P83AG3OngJsshgWkf2vDoIAoH6oyHeIbXMstA4JssF3+fFMHkZvQlQwN8bgYgu
bQABce/8aSk9w7j4BVWd8W3cCanjRK9CXWm2Y59iSaZzhzdkwCfPA7bkliz0UxOr
76vlCgcq9HBqMqvsSVJj55hz3VJIrVT2o9a6gL2EaJXhpm1Kv6blJFDueltDiRjU
YEd3xslQcK4HIf/33d7cV69YtWsyWvnDhpfmLeFbrphnCUmkXgYsb5A8Bz+otzvY
bAKk3RTSGE8x2dVWa1wsWUpdVLHoqFjjwbHKojxR00htDy1chbPOidExOjzmm0FP
ZEVaqU837q8cFQX7B8y3j5C6ehnVCTu+1XdnNAkrMYwCvlGZolGr0mutjssd+wRa
Bi8Lg08V+nokKEUa1eIj4+MkHSXefPG5BhGWoiDKyGMMGbra6Sm8zop3vQ9b4j6o
8FYUXkNGPYxkAmjQnEIDyIv63P3j2by0JyAj3/vR/gXLspkKvqQNpkne2fYBiBy/
KZX8t2PbUTBS1r42954f1y+QrnGs0ftYyoXM5RTeHxH7EBULo4MysZvL9U2XKZYJ
fBiJJGFsnk/TDB5c7Uazaq3DzUkuCFjagIvhZp8e1gno/UghNWBEpZaO2m6jrzbz
EdPi+VcQhXhzYD6LYvrVus8jkRmBzXNARVLyJpXguBQxo5Iwq3iL9g+9Wn9qAjYh
X3Y5LvmfyAQHQgbRBYDZc6T3KQYss5WpDmQ4UnbvnPaa8rzE4KeVTXsgD9gyaZ/7
efYLD7ZnqFdHvZMROEPNXDmF8bWTOj/dt3uy7wCxWl3U5d/m9OZn2PhkLvpslvVo
Z/SiD/EalEhb4lA+j/t2vbWPtXp85U4UBWmplUNryQRU9oEO/odDWO9bXhouzfVS
9QOyBeRjd4WKJiLsCRBoUPkC2xVPyN3Jx8+C3tm+SKFSu/Co6s+UrKGQcdxQ7W6V
qjVTr5HebYtHzC1dfuWTvmSR/B8gjhwiT28yS5v9gKsEZeoVoqS/86N+GMO7uGTH
dhfN5oK/x4YsPwNfle5981fR1UTOKsmRb+Cqm09CaWdO0WN9ZstmP2/5B3b8r1nM
0ZDML5gjgkY/Tm0lRwe91qwrGGM1EB9zmM86dWzpO0NVBgJPl6g9aH4v3P02UMlX
jyw0Q9tha8LiKadtoqtRC3dIcW7B0QytkQIfNFPkEf1jXlzAujzNTSiymvKrJ9Fi
rl7FORmWwuU6dtpMowAg75vfk7KfVeseIBQEC6+LjsCo/RTweY79iWWWh/e4eUgb
IgcAqC0rsFzfLIkzQBXytoM8KJs7EKyX2FMpVWpZyNXaH/mrRt/ogyx/g+3Q0XVO
bmR6mdh3tYyn6y2iR8MNi7RpGkIhMdxz8WXq7IZQpXhQQ53JhCd8GXg5tXETWhaV
B8n3S23w6hBU8MFaB6+DgI8A/tu/DkqMaEZHtw+Iouuf2+D2DRMvLu6WvjptBEDZ
XdtnMBexH5xpiEPSftGeTckdIuA7MWXM98LnDO0KHu3m5I2mWTHFcEkkC8fJqMEr
R6VPH0oMmD8JgOfHral/KIolwAJj7shDRvAa/ZSiL50qX5xf/qtqrEwyoA+vmw9L
whaIAPjTb8E1WGb/lFc5YwTL3nbT1BYN8hJ82CI/bLjcTB3CFwOIcW64Hj3REil2
2AfzUGkecf1gGmfJS/XWwLciqojP4l9scFOHIEpb5vIwzBSEOlQCMuYx+1VW2APV
q2KcYH8qsG7bY3SSDewFogXhddLWYESpECZzsE/xvhl60L4XEctOSgLMnxoIDI2D
/ZBMYExeDbBVTn5e4+yY1C11OOSa7cLLX5WZaeXU1AhIpDsxh/aM2ASPnHndWXo9
GYOoUPrdCzTZZja9Et1/CoyyJVGFAMnJ3IhA8R1+kZJmFacbwX2QBCNoKX7R2AEF
7jpTGc1veV1REl18XAB+KWoQykh77ACFQKw9woePTAO1c9hVURVOZer/3YIIVCMz
GMU++gMGBCrfRBl2P0iXKH0qNySVqZXzICotZZpVYEwe1i/OHWBQFXXbn7iL1NLa
pwwMUkKUVkICu0OBDOp6ROB768qY4vT4Ar+qxWY3hRGevM3z9bYgZGGzP45Bk0Ou
tvvdyP3uoaNy6c4FLsKCBM/kbXgzzcOy60iDRHVkAW9v4gzz17lAmdAGIK5prKD1
9sNJFcFt1ncnufncbtI+qXDR8GI+3WVjebwXZkqrFeJlv2ooBn3QjtT2Qln1AW68
DMjv22LllbODm/EVhWt72gsd0vGPSfF8E0HHPbujW0xrOnrKHkMXskE6+NvkOQiB
9lxg8epxMxl7w6snQy5uBP6SpW6KNWmmuSWR1W9eP0xnLjA0KJlsg66a0ZN6FdqU
qmToPSc2IgauDQocKCcxnUDSE0KXzvXFRBBA7++3/eAyV3FSWMbeYpyWvo49Q4cY
ODKujOpgNxTHT1pq5CG6BaQrghJ1iUywqY5RzuPrvfw53a5KEbYpqEGtdRvNduOt
8LxDNS/rBf25Dw42XiTEumcDzalnMViBWkj7JeLAdIvh8TrKJN+zfthAZtKOQCl3
jauh+ILMVejhfdWf/WWiGe2iyqq1dXozMReBQeoTTEPk5/K4Ilv94riYnHZ6TtnP
i0gGG1WM00jpDCnCWdcJ9qn4Dg8P+jHfPf8/WyDx88ivRK4E0yTIT8neJvn6dtvZ
kRXgy1M3BoALCyUywDyrP86g6jx2B/uTdb/urveTh3mpmtJTkloj6Y8FjkCV04ZK
3J1NNiocFWENwyD2wrjub4wQ0R7Pl3DTNmTj4Fa9/BlGjSGEULgjjquSA6pjObT+
4F+e82qQ5OJ9U80hoSeRsooq5VkXyetSiNSWIRgrUb8tvRgodkoG4nrZmKC0DZLV
7rBl12bjygzIkB5LShy8EPQo+d/pETf5KQ5l13B6alU6zjfv2W+P2+lnjDrYnFVd
NLcsgkTPzI9g91kVK9w7k/ral//vJTCc1bhQPWu0i1qwye84faDz4WuQocmiBruw
P4FtGnMjXQLwgmACJB9FxkWjQ9hzahB+NNQF2nC/rCL/niAhGO7lNcM4R2mvqQtF
D25Oq+n0xkBJl/Hiw/lspUUORkc9qPqp10gWiUZAAAqxqUwYlJ9hx+j818qBEw4F
in8HXek65BZNHKnlQWG8j1A6KiBqbi414XM8F5bob3pR+5X+m+opxfpcrsziCgp0
j6viUsAfewRq8ARoXMb5QSjBKPMRJjTd64sYQgy/YFBB5an9+AzT8jYAHkHld2eS
ww6bgYdt/awbZlpg2AlryQPEdImV8cBaUgbpqN5YON9/wXZbJqmho9ByByPb+04w
aYSuTg/kNj3PjdAtEywFPGT6PeM3I+8SpevZne6cluukgc0U+3xNXQMV7cFhu2AU
5//Iz47ktKSG+yJQZcfJ7BmX4lV6k6Q6DxSUbDYFkHE1wrVl8kAUigg0loScEzak
rbhLg1pgNDrwrtLgYp4FzAX6139YaL7Kl41bY7aUJkTDaP2JK5wJKp73CWFmXrHA
3J2VwsMKJ6zqUaRsEtOnV17VmB4NCn+yJ8sqvqtauAWX48FoYRWIHwcNouSMG8eo
C++UvZf5Atv0zYWKTWnviVR1eR1g+2Y+GiECTFW1uSw1IJ8ucg2j3Cw1d/I6byDB
WONBCIv3dgCvzEzD4g9wpLRSYlZ602sjtftGW5aDN5oTkk8MJRbAN1rVDzzz7oh7
Dd1x/z9VhwitLhH1dgI88n3hULq5VfHUDoAXQhNH8+wAJDgnvyvuliU1mUBeGuvO
fuSLII9VozL234JE3opjekpz2p5a9Jy82UNKgN3itw27vl2x5AZG8tK5ZeuYeVTf
5f1FuasZh9ZlV6qv3jW+Q4zSAAQoLA1/lC/0Kzf9UWENtSW+bkHD5A9n1wgHff53
p+fvHaYqNmZrSgPeLeiGnCa8bXls/JxBKvzhW9PxWHXmGwagYL00/LvR6/4QPCou
Fpzam4JQRmJRc5ljgsQIKlGEstCByTurCh0wRGr5sIHHi4SHHwHnRP2OIi9A3hII
/9X8MQElcDqUvE+6LLnZddO6LnTNlR41X+UKUlTuykHqKxw57ka/lVfZssrHcvM4
gFsoVDuHQpSpAKPk7Hzfd0ZVNZjSgqZ6C9hFAbzoivLf36eMN4LFt5tzQQZKGUok
NCs2oGArX6n7E4+01zDkhX9XEVdEFBX3O+y4+m10SzDjOS4sLJP4rQAkQ4qCLKTz
/iQ7bSWVaipOidz1UaeMy+cEKsVdFLNt9wVwkGbXxHn9UWMNhMthErO6uNrvYHv/
qQfGZa4l4mLTciTteQhAXnZDZHllavFAjp4DvERGyycgdGHw3w2OBcUCBL6Fy/td
Xv+6Lu7K+5xu5E2jLVMGidlvIo1ik91qhYGIYVJUWYaq1Bzt+aBNDMtHm5rYzUQL
p8jDEA9m1Sej2N5R9xlBs3xZyuOLkp0sDqRDCnIPRvusnJsuoZv+ydQsZ/UKXxaQ
nzY8QmjLz6dsBAIyZyQLQctNlxtO+o5y6eyRoP2Jlt3OyqjND/fA4zqONXfmY2DC
PttnSGyJVc4K3lxx3cFasXtpURJi2ivU12MF6SxpmKCHEtYSNEXcvShkH6M8iGGm
dc8sEUxuB4m/EjVM+gN7pCdLXgTNLw6IK9zzDA3MVMf51YTlpXybXfRFtKIrlL/Q
SG49ugpIRgTfbaoKYN2Lk+vCRYADzRS/hgry/6j8cjHzwpoGl5qh+drUgNOnHwHU
j1otxFTXQGPs+IZrlBvysbtNs8VX+oekAh5Y2u8rt/vDnGe3+zDNsUNPdtnKmfE/
7omLj+Bsh40+9iAfTR1dFw==
`pragma protect end_protected
