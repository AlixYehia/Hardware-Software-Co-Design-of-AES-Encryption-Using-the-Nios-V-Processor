// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tULFgRZqmbtTr5RqSVjz0SnLGQ7eWZvTbEKcxKhRPB/gVQSda01BFTrEUpNaItNWUlxDe11sdVWB
MMPOYMt4pb1hgXNAlzegGa9HU7TK4Dw0Dwy0gCUepfmccTakLTAX7/kVnV7yrQVR10eSOd2yEKLg
IQhityBiG/L49z817qNOVgSvl6ppgi5aV1r7/NmB20wKPdcOhtYG7J5BpXvH6rhxbILk1OWw7DYt
3NV1pet6mQpLEw1VLuWZqB83Teu5zT8YI9HB2BKXW8afaii+G2Zv//YylMLIEoNVZr2sfGI9NSo6
COsGKx3o89IiTpZxZZ9QXF/ZVm4tWtgmdcd1ng==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5136)
aKVG34D0V6MOeRQbCz9K3gc4uh1ErpolUvlvg26/3SbZisod6KtVuFAtWlAdUuj84MfFGBcBmp7t
0csz18WyatBuYGUFIK+8z5qKR0g5v8xIXUwgTOqC2bGxv42xbL+C1EcouPU2blMEnxcSbzspiN/R
+H1DWU5fQZ6RyoUQatUbd+3glpvWcceqAyP88j4MO88CKRdfxBYANbgS98HMlddis9CRpIgu+XgK
xInAHa0Yq7Lkz8urPBScL6r5jOfLq3eZzYegUHHb7NvmSc2raIwpiOaWb4IdWbKoKJAlDIuvnKM1
q7PiOWUulBHT5q7TwDDxfMgF24T8i6KmM6ffjOH3xg+HpVX5UpGtkoktda6jUNAxdRwYFftFK1k+
+K15CgEd9zAJqp+AroA9sfRZ0nlb2pWfCxyOGQNbvolh/Lu6V+BC7S0fUXpC50RzvGsvXJWw91hf
bBH8Kxrwx09xqMXb5m490Ys7zKO3FhmC7sLcYiy6KTNGe8MaqwSbK9s9SHqO5A3yTSujvlp+6GuL
vsnFnxhvK55f7LGRNwt5E0RYDRXcg09hBiSNAEtuCLd4lIx0G478wY+WubSXgwdTZ9PKTbZ3mmBG
oKU3N7sU2RIpE6oaAy3cMALjhe2m3eKupzbTkBHZevPT8IjENrHDmH7n/x3rMZWgvAkSGUtbgBAq
W3i5Qb8O5UsoDJMEpsrb+sfSKYMzEUI3GG0yufE31WXC+ceGKyXbG1Glvesrx6hSEyAVrq4gZ+4w
ObMH9+VXBQ+jWEx0vS7R9anR02waLCWxiz9wZvJpByvZfg4H98DTW6pLXYzbvYTmeBC/QHbeED7h
YJhbVTTwL/Og6a5C2AtgFgGC4CaHPO5h7ZzbsnOYqeu5MeXtv0IW5zkBMLiYoNnhDXIoPQ/dD1S/
mDMr3/LQxg/eiJGlexVMAzn7C8PSPCN6CBlsZvpwrO5CS+iWCdS2VXl/dLe0RSjUEAI+lg9n5Z0R
B0KnpZZNzVs/9ngptWG6rv9Yt/mP9BHvFKq8O7mxsprLmVf6cXQsRXhc12jS5J/OchnNMvlR+jMk
xqCGd19T+nxjVmXuz2zvUIjqChjWcFfl18xYQwUXx+tzr6ixGz79fkRIMP8JDGRMDuiq/khF0YO9
kN2794xLouUJv8AHO2mlKCaBkfigh3E3i++PDtx6qiHA9Hf5eI5bPfC3T8+zfDUJM9E4AAaSHXVd
6f97KztVYV3FFqvnBHpSCTf13DxT05IT1sp0NnLBCQBOWYrAx3uzs9MmJXk/ZxjmNgO82GhnkMrK
fDXXApBItencuJQNd0UUHUsezNHm3i3nT4wpYWSOkquHzpPGJX+fIZC5Q/j7gvsNFBNPzPuH5w1n
6hzDUs6HlRqT3lRfo7D2d9DQxos9Covse7sgmThU8HLLaRwJuyZowtGPfj3wXCW9RHroiliCpyD5
BDq+iW1nVo7nv++EVDS7TJrypAxZGpPNyxsLsIL/qODDdXqPNRIG1VxFsXLqQDSSbR8Y97/yxy/D
vv95KTsy5y6psl1C9jVeoShxESPlNLhmo6u15BBf93A8iLdYtHK4vwR2rE0AMK4GJ1Bu5AZbbzwd
w3ZkS+JR45ZRRj84jR+uHSfGYQPKLJFDFT0ID1aT51Qy6c8kkg/V8ux+LQrfSqv1LRlpEtb7LrvT
5JhCrVXBiCZv8uxw7ve409lT0Q0KHDtTGaE596xQAePUPKejvuhwArpiNF1w6aEWByhpRpDxiCiz
UPqExvPO3efCklT+DuaWyrOpeZiFE1nnpHkTvsn42Ej7CNg5Z6kHHkN8ZyQkdbPtL1XSs3Ij3J2I
ulY6vZ55GgMfmM/i/48f0NUszFF0yNTnw+x9zaq7tcMJXgWyrUxnYbpSCN1aYFVO9AEHXCmCDak6
K5SBBUbGEbNQT3VGDE61s3RgW3NbHT1/78EwJqJInzrmgmBhCdEMGOW20zhAZCptjzw6SFlFoJk3
ibYF1he+nWDn0Fhoh0YTWHaGJic0n7zN7nE6zOsBwlVxdoHks4nr0dzeHBIgQ4GIBKRvqYUo/+0b
3ocZE6GJQXJkkq0X1scMEWNkEpymGGPfGpaA0jiBoyd9gdcNS1kcK4RKiWRNbU5btkVgzWijVEua
RFvgAGof9Ub4iSJ1npt9MmimhrYM7C+H/O2GKpwIi77QMxrULR1c0VQ9AAYXVewLavpJoE/xebiO
TyJ6+z4mzwt/I81kTOuk1u51pTrBSpCS9vysb73c4aQAQkUMj2kvJZTd7N2LvdCYMyoN0h5uhdVW
fOlbl3PCqslm2p8etMxYPZAhLj9G90JjDhKyYboSFVXnQYXVoOEeTS4S7wXIueVkdiWh/iipkAtn
7Z+yAf8Y8eueddFUyHYqOKa7Bm7GLRUYngRRZRFv0MXZHIVM0DcqqDBT8P5PAoNNtaK1tJBNSTA2
jl67yq7hPL9ZQHK0uzqpK3Q2XFHUefFfPiY2LDJw/UkFLpiNFoDwmzyHBJNU00U3gI5lfAkcjeJy
xkncywOuXAObrfmzEqb+t00KuIUGnMgUuB6lqpKnZeD5wYIFifW3W/p7spJHHYxKweDfb6B4vnsv
p9D3tJsf1irnNphwtv3GGoxSMajLTFvluWpdy7oVbrLBzaJPkP0PhMPE7OzjeZsQFPQlAURC59H+
Chi9rMvkRIBkjbWIucmQSNWskghlo6emaWO5g8OCGft1vuw6OTsDeTo7ojmw4ujfmocAClU7/zJH
/95LpZEWgCVDBNcqtu5j1GOrkIDAr+3TDPxBY2uxGajZaHgxsRJdsxP9UA/VKQ2SbTvzF6gTJbdo
A8YU9Hjcvq82enTSmwqoRFD6Kc1Qc6LP7lf+jnSgs4zTEOyNuxmJddNMRuqniT6ZrGFUJmBthjld
NPTZGQj7+IK1Lzpz6QCLMrMbaGsmMvj87sk8nNttS+FV638EkkWYlTdDeQCLDTr+kQbEwv1aO7uG
JgWg9GLgvOWDDLpT3RgfWZT7VG+zPRqrExVXjtvdnv68dJ1+PtNpB+FOYI465waVw9w3YmU7KjXE
hyfkfAjfyqdnF+yqcge/Eb9OymM6qLEbTQHQRvhij3orXgu+eSgYiBBYc0GJ4HhF0iouUXHPed/X
Jwn2JoE9UJrTQb6ALO0GVtRzcNP+7oJn9pC8U4DbIgah6v4z+QDtoSdFhSQVEUcjRmEB9mNycpIB
3/uDhq6U5653V0RBfcyHuQA0SF0Ed0yDeZytAMeQT+pQlrDdFoesMo8Ch7a4DglvjGRBJV///5Xj
BNoLKslx+t5zbZ3jXh8f0YT5GHq/VG/hNr5WY5pBh6yq3/BoT417O8+asAREYbAHi4tV7Bts/MKs
GkAqS7U0pdS9BP9LwcZnRDq2WVvSBI/kUxvQM45WxHsNBdNZ6i8ta1ua7EMDXOSiwdfLpOp1lbGb
eGnwIhwSF45v52VOgRWlN8CvbeLH/jq2aYw0MRlNCZtL/DOYeBYvmZi/HiWSj/FOIjhVJnk+GAXk
s4TBqTQbU/XrcJJou7Bkou1atW9/9XEo7kLQB+cs8T4QsqaF8luXp3Umnb5ycqe02uKe/9/+kyKa
Xurz/FuqWLUBR+vfntuZ2bj1QY/zOkmCfWpTxHIeEMQhrXjAIoCl/32y2S4lvUu0eJhhyjht7aoC
95Mmg9VC3Ol2bGmHtg26pilEtFx92dRX+/ScGxunX1Rgi8sYtQHh+/lhHfHQOPx17UrlUxXiCxUU
6ay9dHgYl/GGRcRi4v/mrnH+LufnJzMnP/2Ph2Z9bgbdrGmGmRTy3VAAmT86jSe0sEmDmTnlpWRi
1s8uYt7JPlxLexP4WkkGfD+8wj0eMU4G3OqciAJgz3IyJJgmIlt1dQtoXWatSGmPe/EvS7oFNjc4
+bchyBU3CYOb+CE8eJQMp2UF4ML8zK27Ta9ic21I11qECZwP71c1RIBz283Bc0XW0CmUrLHec3yf
t8GDp3JfhVn3lxLQFWVKpcDhgzv/B8CqMmvNPYYg1gkTV7zwDl0TxS3Ss9K55SKO5vA/ZpwyM8ic
SXs9ggC2LPF1D02zO0t94Ab5Fe+q/VG29YDup7DChBss9lBpVvd6HaDjEm9IyVoPJfxeWmndgBtS
fKX9gxm+TqC2hWyZya3vdHPZUzoouhyyi1gCoUsUTvquoWU9jiZ8OM60ATaRXioe4rU49wBTKWSR
x4p1t7xvu6lYeK1r/ZpVd1d3ex/TVUlROSJBa2H1kyqtA+LjCm2KUL/D9tO12Sapctp95viJNcZ/
kNykzqOqUQFD+tiVzByFdhu5GY3FtoWQt3e4YQvLp/O7l1JJb3F2pxvti0mLSvKI2VSRnzDKWngm
SokznoweCU40Zkz6quIxp17H1huC84F0m0AfLz/hKXBhPQHCm33FYimpwOquC8s6sBc50GGYI6o6
clF5+GP/DNcvY21DjqhMVH/WWGvKEL+BKUFUkm90v7I+8FnqAIGkovQmUMxWOieJOlaw0VOQA1Yt
Z7GbfeM8As4Ub0e9McfQEaPIZ1MIlVMPXn2S+RDd2JMQmZes3NfUPKXwNp9jz7NOJe8FTmEW4vVe
Z3EhP/DklpVMtLBnIV/DYC9AiNwHaB0IpfsqBIFzwpsVTO9NVcKcuBrYlmFhBnByci7J39Wyv9yZ
iW7flSUvW6/DPo0DyiDG7cYZNYkp4f/cSW9QVwOzf9ZOTrxHBl5cPrIhJYGTkvY6zGFXTOcmCyEV
4ohdrUkJNSMopCEUoM8G48t+mG33ngfIrOMG3rXWTDWDBiiGr4XEc04wlLcQ2gGrFwmuUDmd26B7
O4sIpsvaES5xwbTv7ddLcb6qwCz8BjP1w37lLKCGa3QxKQ+xaUDZ8odAspghHSeJL23aR16yh6XX
AK1LpV8FsCV9rlU8Kb8hxDUGizFaN0A6NrUYoo4X5KzMGNBp+S3t1nqIZv6Z1tPI1TKyot6WMVqp
rKBQhESffkwDwx1DC+sK40omw2TCH9h3kAEjf5dFPgU+jQgONgA1GKrdvfJg161EnkKU4Jz0n5Jz
9XwgZhaeEJexsscFUeUuEs76/Xq9s3ooQTNZ6XzObIbTmqRuKNhRF/WvkDEHFdlvs+rUw22OXxpY
y0H9Z7eIylxiPslstQZp00pr8zjC2Al6spSsrSOgHVrg03X+QFNy0t1o4mLa2Mr45Bx+iHkXS7ht
XM6V729dRNd1/FM+paFAgt4hPfg0Rm7I4RgbxY2nqMBjnGBjfikadWQgRH3L9CvKh4mMNqELAG1W
I4xGzNTZ1mV+cDtb9+l9CCRkf79ItjXbYwnJYaM5T4xjWiP0QsIzC9d3OhkpZLq6vbUdMekUm9K7
UbluRTn/ci+sm6MCy4ApI/AfSNU95bjEeRJbKb/5eSTz+SeGiZqxyBKfQZZcIRM3ZW5BWWdE4L8p
wXpzw9Szq1RW8SEJgEDXAhyDAo3g78aAim69dxh6ZKQxjC5agWmRsYZQ60QIylHJ3CyMX6A9KKXb
CpucxZUuSfO91zuktgYFXIzeC+TVR76Q9Tmzk/WSt59DK7mu20emLdgVR1o7I2KXM3AeIZJ9/6Yg
ccpCPnmP+/EauFmrM5pLKTqlQMTFkarUV8gmjIKmF1O5eA9FK8k+vnxjTXzueWVcI+eBszE6KLkQ
8K5vbiP/Dj7tXng6tinpg8NuYbQhEGnKndOmouKRE1Lj+7zxdcJdGIfev8lbQ0Wpc8fzEjyJv6dQ
xzejQcaonDsl45BZF50avrPm7UXUPQfQGAxnMmxj9ZaIyuwp7yOe9a3Jx9OUFvt90wFhbvSKHcFK
LEfnAL/rCdFYQuiANvEI4Zq89yNwohlW3U7unGhcZrh2+axLpsOqPwyOVW+4j7dXsIRW7I2VlJ6m
KJlrhdA6Z/hIhJJ3+q1FOYlpq1Lgu0C513HNUYHzcCKbBGIgt8UZrYCflBoehAakzdATFb+kb/WA
onAcblJSuVSNAHVrqI3ZBcRgSp5fqddTVcJ7PbjWEVfhNfU+6a+0iahxY8Zp1+hoYbpVjzalCmNA
Jl4KGjGOQ3jdagzU9A4zixy8MdPpuGe+7Zbe1/JaJKoqBpaYLxj4WG8lo4l8tGmx+6n03blxcXkO
6wmR2pLdPkeAwS1WAwlxvKCq3aCjJXFOBUiBBFJ4CWoMYaMn2boZD7NwLCMzwKtVRbIEpq2QNyMv
PmmPW4zGTJKTwGMiOdiQwQ21tVc2nuCxf1TfHtEs678s8/RqfSIhPFZZlpE8/wekeH0diglHNOQZ
rMXDERYvAopBQX0IVnUQCKF2EW8FCmv6iTmOfc/WP3U5CS083SZomPLKUFwZFhCQ+tmLmmyyGVMy
goRhwY3NGoqM7oekvBgl2w2r+43CcolC5dX+eoJiG3p+eM2Ed9tUCj5VEe5dEjHvYsJw/Hns4aGC
qKAcGjHCex8Lp+g+JYcbcKhmzBzDtozxLZK8yEf7BCxSR3ha0mH666wEaDdLBcAUlsN+FCFS0VzO
QRpBYZmFnpHBbN50iYHKKDBDYQVMqf7ZZ8b9+ncMunectesyTJEsqJkd3w8DSJHyZNrgFWi/TSdy
yeKr+Rq7hz46yGl99Le1JMh3WkbmPRt3Y8vvRyUyrdwubebEkG3/WzVuL6oAsE/aa1O2SHCgMikW
miOugESfmaOOvxpxvv2r0BBpJo2TI6SmqyCbL/1J7eubvgdb9iv7cCDOctrkrKBaWSNK5PwmxxPs
5u6/Hpoi686U4tWwPuufHTL/PlWEVzsM1cQqmNO4bK5/zHPf3WoFbA+RCQGbAfZqSIivcuXL7Lpp
wWNuNdtNRveWFi4g9ktavUKBvShINX/2Tv7JQRQGIL7v6MskbmIPXmWEsccYydkUzcwdboJMQNBH
Yw2/eE5P
`pragma protect end_protected
