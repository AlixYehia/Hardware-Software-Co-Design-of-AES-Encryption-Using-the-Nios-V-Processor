// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Kfo1VMTbWzKr//sPnDwG4tKb/JjMP45q9S0uxeZnmMzMBX49YW9iHrraHT6k/4P/+iw36CwyUss6
9RlImlRIgijz16/tAH/MSmWrEKIo3ylekVR7GKVhCHa3FLrT4s4UOu7jls8A458R4qb5FJaJIRRt
YtCRMkAvN07RH+eZCRF2NX/KvmS9eD7WmjnFZ6AWJBuMQv4g/XsbPskfjFRI7/wUIfpunVgRUkw+
frhyd35EH1S8so26CSt47sGfIsyumXpvE+CktxPTnQ1LxUBHmceyfXam40XuNnbg+jOqZ4zezn3F
mdPXtM6WxYR7VPTZVxo69XrJl/kprIMKXY99jw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15552)
oTQ7fAothfSPHHKqRHbe1mj6RUWDolbQPIC16/W9IG/drqmbSY7Fz/XATopO89chaXuHRCpNkwEU
q2Eb2hKWuP5FqQ2K/oUiuWBsCZc+KQfJSIhmx3OQVM9W7kUHPfUGChjxRpI0C6pVuJHBdtzmzQdz
VoFCPkoSoQ3jXcW807/WfnXTTtwxSP4a8ZYqrm0KGbadv/3EsP3yMRjPukdjNr/PSlhCZypFDKqo
dPcxzOFD88Kmseu5FTd3eT9IqbIvCIIaM+zdzPr+8C9jxIt5b9sjK4wYcZoyI/sctron82f92oXH
TDmSJqhlDbNob83T2fV0EP5a/wQttM/P/mF8dLHozvctawgzTz1Hdj7qDF9y+v2xX8Xr2aYuF4jc
s8KxFIsHTnIFccQ2tRY/hKTomIuubr7cKVneg60gSChI1oDc3msULEggO8ouc9CfxCqeNcwkGo79
2VVDzW+5sAi3vdn5vjg1XxFYBxz27bwAL0u9yXsyl95/ZbXejydvDZa/MSM+dMg8zeggSWQTOjq1
PDcdE3RL0ZgZTsGk5Fo5RgB8kys6ORyB/KBkc5+RqE3m/0MrHmHP8LdTPGtTTGpzvKafR9b9D68E
E+FmMKlQCaAKfiHVVegCDjVAGpbIY8VeVvn/9XRxlc9sv3vVG3C8A68LGMHIjxembQ3xbqoyLFlg
tiT6tt1+WCL1TeW71Ot4ZeQup3z8oOHxknhTt10g8wAoexiA05fUbwhDVkHOIQWrxjZka9fzLv/5
ej1c1IgjQ7B7TWv3LZnw7nJS8EVFKWiCp4Fl1GsZzPafqvyJKvrJXgbCzbWu9BK0xF8+QYzFfRt0
ua7WYTw8gOc+Znfb8rXJaonnaNR9Y0fixStvMe4Zrr9yA/peWp3KQhIW6Ve3lmCHVXAtTzgEfVS2
mRiIPABrjqKksO35ZFj510LM30KdKGZ9F9hy47bPlEdxbwfxcpOldMIP6oFeZkoxxY0x3pQLJ6KE
RfQ3lOZc1YGh3r/phWWZGEZnv51xbYLrRSMmi4oS0pxgDJg7N7iCp6YIXn04VjD3rj8GAUV65xt4
3lxE8tMmCLanfUVkpLSCXQwsBT5QsS76sUWCxboGRNrVXJfUhRLdLK+96eacyA3uC9cbe6o9US2l
HkMcq0MMRfdwfm8S3/dkRznDM6/9W5vpVVpB9rur3mWnWl48keyb0uixNv5yRrlVBJoPHB+QRO6+
KQV64mQjsMysJ3xbC4iQfeMQhN0rk+gArN0XL7bv3SVcmJyGWvWNJrGtcUWDKF7AnNZu0xIOLhnE
G/Gjh5SZOzEyqhbE8GhmZMFGSX+jpPQtMODSn81235fGRl5y+HoCIRk3H0FRgTelpamUkq0vFbtF
7cenIioUZXJjmua/3HRQ1E+hNyDQZeOV364FtLCrVq3QigDIxzOyBR1djppxeammQKEXf/gYQp2m
JZaYc2TM7prjGZPb17zDbAx13x1248QFJnCBLa9xr+F/BHXQ8nEhO0OCCDnKYkBiHSdF9PorNPTY
Mo7JfsRdJ80Sw2ElxTbxEChymRkb475H3hkmSmkPhjYIHUVIpm7TSu9Dbu6Ofd7unekSXP8KdTpC
ipVsFuVgCiA+Nzw7NdbOcoTlw1U8L6RiH8PI/mQvBu/muMDrl+rV6KeluIT0xoS/DfZpZQ3DCWYU
woruBqllDUGgwyxvlC2iS9Hm/xDaPaKh+Z3o/Uhu4FpOBiekA0yp50X8d/CeTR+km94jWtFETTnU
5cm6wzq3YaQHPRgzmiPDlK54g6EnM0hCijQ/CjKkv/GK5Qf471h1/fP25iUKEk3Zb++jR6MYHbL0
zwo3+8nxEszfEp1RrtvgLqtZ33YIrmRBzixQ9eX11P97GqSMZzsR5ro9zuXUOH2T2/1YU7wXQIlA
E6dU0cI4tLpuYnuwf5t24XuFuFcjq2mdn2zH7DB8pWn3AJBsKLW4G47DAcE5bCQra4bbBV1J08Q+
0QS3ZWsEiTOaHMOx65kF7dXyIJTe5ckROsG+/fnya/Tu5fFZorQWYJr/eRl/P0THNuu7mKWziTSX
+OdyviKY7NQlvbsKtMXq3SpwE2rPfXir7CAV42YS8t62S6rBfgpQwLnU8ywiviBd21CyzoI++tkG
paSoV5ji2VNgBaPRJGrTmpnVvVDB0Wg1cGgoecmI5cHLvpwOIqZU13U0leOIWG1ae1Z01fTkpZXG
t4hBWgm383CY+QgR88rID2x0XORXGFbmMiMH98s0u+7Tg/eonGhpw/SgD3D56roQ5eYG/qHKpeHE
2YWXDWmclSyNSOSGQH6/kro+9BlgP3u87c5ok/bBtCPqc5bNn1fOs5/mmNe5UXO6ex3aOGOcLXnX
EwCCTaE0MJh4Y57kMnYTG5UXcNsZa+VqH3msT06BM5G3IDhBlXE0dAJwoKlRYwm09IcdeAeqxvs2
fPwy/9vgZmtJ38PGj7ww/7AiEJZ+r/ua1aPiCNHMgSnIGl7w7R7DtamTYqX+w1/7zhKKSXiMh4cD
/p50MocK53L27nyHzHP4lzJlgm8DRupCPxQGrKbfWWnhgyL1jtWE8r2YJU+6FOalDwGuFnScKv05
Znz4BjlAPzJPwYSQa5Eehwf4ZzZJeKxCZn6PKlsHMlyL8X/cXf5nYB4/n/bxUG3F+GnV5UW5lotx
ohwY2s7nHDOQieFXuLklv51KznfuAqKBaKEtkCYMw75mflHQCWuh/hHcfdPS/TAkYi2Hnp+ukwAg
7nP+OM6zPc2tpTVUm3t/AGsXwZgWWNf1ozcPUuWxb0nfnPZIPU8QxC5PEvKZ77H5Y9AXwoR1b6fE
LFdMLZzcK2RUb/vpOlJeodU5sSHtvvKeL38wnS9dKY+ZK1jovOLJLOK6xsSUJwajxuZY5SchqXf1
nheTPk0pI9Q1Ce9QAqPKC3osskQgFQyuehgAAErakiriDuX+XTQC8NkRpd4z2HNSko8YUOOpm8C0
yFXOysp74b41GXHYHuEBDIXdqA/oORR33QAv/YX91W5NfTUYUe43mkWeV0Piswa1YlTOC/2M6rKa
J+mlWeXbu0TTb5FOLK6kiiVmiNr7pIo2Fr9FLVdsmIXgGmURjzSwgZuj7nVxlsP+jplKcwmyH3Ab
6mA5Kzk+xgwmZhNlHPut4k/NTp4GsXpOrWwAKCoG2WPITXi6m4KYP+pE2i4ESEkvmseFSOf8is5j
84ScXqNUBEMrNij7O/pLyRdv/nEc64laOov3NJwAn+kh7CmjYlqAk9cEwPiskY3pxpJVKkSNx6B6
ah8QvWupU5oyMukPTBIYSg09HaxaaUbLggL+7UrbLXqJPNwDS/2rfG7+VZbTPK7kpMj2a4w9vRjS
q+gSazJk6D/f1VNYsYHAyNQmsNU19gLI4Mf5rCV+8osby3NatzM+wt8rhH4KIqfKtK7XlwjyVTfD
FSki9qiERx1x41cNLVZEK2ALf654RAeC18DZrOeS2uU1vziBnTGUCoH488web3GzrC7jK9fP2c0Q
cISki7aATvG/qrChzin/bMu5GAb304N5GPl5XnLx2vM2OENu5NMekZuVpRbrlrDDceKMiqsSgahz
u6r6Skl9UbpUoaeftBUmefDMj8EaILRZdmtaurlbbBZ2igJX5/4nZdmktjPMbGhZtn5eWB71KPtO
7o43TmX9rURzMAF142AKgCZ3na2AyqD/b5R99ZpYMwOa5s0xIrdq6b5VHgqL6vMoLjJ0VS94xknC
dep9GPnukghl86qv3KsK94PYE1M8vsNKr5kIJhsHF5euwOMEQImTS66vHi7l565hQewgWzI47eUp
MI3oZ4hqxtafbGDNUDt0P67R347GdjGoOEqRgiMvGLyuYvHjllkudtk+qE8ktJC601gZbCLwPqCz
+mfd40fhgqZTxkfDkIS6DqwDTv6pcmqmP1n4twSqKx/3pUzXn0DHEpmX7m3mo7SwJSeYWC62ug3h
VxraQewJZ67EeSq+OuUzvODHQu5J3Julo9yTn8ghCDCRdRMPnkwkQaO7CaiTiqFVpwGpfsR/M0mP
WbOcyyciilxx6MI2d5xmVA8foOxdtzM4g/5nprQFaoRFhT8cAgDDezTHNfkF7qb+Lw3cIknteZsQ
qmIUMeDxXaXQvgP+B0W1nn3NO1Fegr+A42GfAcUBVsS1A9VhHEKCaMb+y8n3LYKCwq6r2dnCTgbj
c42BewM/iTAJ5z5RFoVP3sX6p1gnWqzDwrZgxlkJd8xKv2lrCPW4hgz4LLMeWYPYxZU4f4ODUHYx
+STjT2qZuCY5q/vpg0Kmv1KKFQEdgDELB6qESlv65GK8iDvpfCaKlhdNGGB60fWf/g9MhY2XpEr4
pehZ6/jn8vw0izQnAfCpstMUFLNITCdO/VS0Q+EVZJklEV+HHP0EniCiXm2FMo20ccYitg3Kvltw
m/Wwx5yLtM9yIYcJZymf5SnJlNLYeLxh2b/sqSG/sWsGKoHx9n/lRODXC3VaZDqcOA3Yf7Z2utVU
pThN663DNI6e59aQORN6dyNu/7lACf8dDmB/MwX2gXflNJm+yKqG0PHthyqaTYysSCCwVORCihz2
S+N/KvxcaEW5NR4otv3NeYrpt3OuO7Ul/8t0siWr4GlNuE1zwlS+nYGb0aQHzEALLFlCszOx6Ic8
FlwjccAJBu/S/of5+iRu5QZxa2iZjFbfAymBMY9eIILwiOprjGsHKX24Ka33rWSWoJuKY9MKkNgv
rwl4wHrZukCpjccIT9JRqoYWGShkmHK4/YrVdOQ+4N/W7WYZWpeZTlko2uWVQiMbibZ7X8AmKj4g
rmBJCfUV5L3B+SWnw3WScixhyRgNLW8Eb5lcc1e6nsfuNdvnNwDw9r8QCZv+Z1Cz/ktW5H15zw/D
DjnwvYbb8HPnVwlfMNFiG2nV0e4S443zIsdNVkb8L09sovd++/kRtEYws/VzwwcBOLRnKNsXfmsS
Bal1oVxVZ6tkI2g1ha2Qt3oqK/JW6M2HHOmeCmIUxfn8MKML+Ch1Ain/gPxuAzWGDpKVP67Qk3cJ
hyZqznVMxlEZqdA8Ad/qj7EuOqgB4vMjWd86ptoW8aYpIDNqOfv5ZitxJ0zZTaUc3HK64t1jdZWg
WTASQDSa9li5xwTeAhvaPAUxPzUIJSihqqvw3Rada5t+WIyXWlAsYTtzl9oPjmu2pp+mal7ISwWP
er+Y+7soQqmzZM8eqyN3lv7Q1eK/2NV1jth8QKCXCAmJafjGjYIPMKptJD8wxZDKl8caUkXdqVtx
jcUY4elmcIulP01usk/LBg2fdSfC0r0vYk2pVEVNtS7pD6l/MXgsDCX4klP+ZnNJ2PVJr9C1O0Au
Ozt6dzceqElNY/FSA2uy2oGQP7UVy8RTgsgxjJefZlLedxRzdhU/QfAdVgwOPp849Vr9Ma1BFghr
raEuyzydPAYJhvi/m+NTcSGMqg8avUwqteHwNs6puhsU8BZkr45ByWkx7P8jqN4NMnku/blADrO5
7EA4IjXO3mwBWJdgl0tZSSrjdWBEKdLDpop3Fe6jY4uAl6TxSkIuK9ItkAAuPSW+y1pSkVyKhnSN
k19GVC/Sa6p4DDTotkjMMEiKZNPD9a6MAF+LJdA2atPHYsR0aWKYObZej2+112JP0251t1MO+PA7
WF5gdqt500Q3CpgmKx0WmO9+9imx6OExMtvMMGgFBCtUC3XF3scuJC6Exoh8OnfIG3XF1icnsWYZ
JAzGa+DPklQ72osT0fk+300iH1H5qRGGxXinE0p9ptC5gSAiXqzQZCCl28J06TXhU3HWiy125MqL
HQHtQiF5u4ec0gK/kwdiaoHFqfp+KTici9mbbFn7btckhe9ZhGReDB2GGAnIm0wm9ACGZHx0ck+2
ypWvyEpSuJx2ssWdEgOmN5+GDOEDGnDDskcJ5jATYx3Tct3uYX8/Hucd08VGzJ1zT8h2y8JkqlNv
Z0x5QOpHRZC3YEt3ixAmGIxGts9iAnicG4s0+qIjKty4a0FNVBCjXUquJkxj42GYXLYgbaSc3CQk
OWyOZrJlcw2NlMKngj+IVcAaxQSm9rL5+4kFja3zpDAeDnKpMSpy3IaXk0ZyQw3Iigs32rezz4G2
xdIcrUkQnutjU5JQjkbWVK84sq91LC6hFQtANh1m/wAswNR0s247oU9oVOb3c+Fs2zA4cUA/wg8e
n3Nf58PkV6OOlaHeciY8a74zrzhrda1cVmCP+vmqlFz5B2hbaYmMorA6XuEhMtFSShcaL9Ev+o/D
uhAUevFWEDmZM+XXY9qlpWzwXX2UPaX+Zm4NBMxLXcnkmiva2GYRsOB4C1wFC7Nu1IjN7CuAktR3
I0Oi9oHa035vb/Mo/TNLFqqqmWe/oDc/3HijrovO6780q6J6vqfQ3q5GLTQMNRPyyVjq8NWe+umh
YaNCXEITHML7XOkd+zeqZNBKZKyD98pWoYEfIcEw+r/uSIJgo8t66iZylWiLiCvX8EgrgMCIZiSz
6o4rOgfrjiW9mxzfWDVFckS7WIY+TnR6m1uYa4OqUcbxs8nV9GqIiZ7a9iiAdsROSt9qCrXrcfh0
wsziG1gefm+WFyKe6YeWhM0vxLnqj5XTFRkCeaACIFlAAfktRMM+JxV6lhm9t2CyJJlVUO7+k/EA
mN8N7dqfWdrRb1hFOucec/SPNWCBLEt2+kobh82nlTkbpD5PfKHHVYi5kfcqhyCVpJJiFFv4c46+
CGcDeRP8mpfoI0+w4eInSlmxYdLvUBWCbsXtbQ97RIoxyHcnzX47MdYCx9I/bN6A42euoSu5cUZn
+44GJj9to/NQ/uzotR8D8e5PUf+oh+ZkZaBYnU3MsyFiif/qdrhC1zqszscM8bzbZSxJ20Z3zXcE
kCiGGWfdlj3lNV4D6LHEBjRt9JmPI6SWDeBXQhrONL9r1bpSm2lzuTjMFmTq1/opu74sOLT7f0s4
nWrzjLUvT1jrHEeU4q9Faonxdo9ODYwSHpKv0UPNJtEDRBrJxyOnIWasfwGT5P+8eKhGxWvoh4OU
3XraK4dWhR8D1rkVVzxOwUnN8yY+J2sr1sRcbXLOfOIGWLu95CzqGwxSxbz2ZXeBmjgPgeNgN2D+
cnn0ON3VQqEmXXfE2sMTgMswOq6y9OihQ/0HwBo0lbeM87azJRB2k+URHF8dn0TMWPh3AtXIw2Q0
nUALN32+D053Coxwwpe5vOnncFKR/X2Jh8XCeRTWAqgkhvM/y8HnYCVhxuZf93ZHZJ9nbVSXEN+8
0oIdXt8Ttii+z3X0szhGB7BTgnG8K/0MVdKg+AadJbAMyen+DIwFWTe5yRT2VU6CjXBZSAwCcIe4
9Pjf2okoJlNk2VirpwqQcc/Zod3u3nDO9YIh5viAc0GlqJXyx121F0WmBsywgRFmzmdk1L5WG7De
t29BaArtONs35OCMIPCv8gSJDd8kJdUeuxKealpu/4bxIJXDAkk1yDCWijHEbTfRPDQvPwNU+4Bd
M2LOWEY09viitciZvcgJoTJuTNbhvA9CvhTwlJEL+h2kqmUOop1otkJeUi4qOdrbgRkiGiVYFGXC
Soks1sQjubVtpT4WIbdJ5XRD3zq4cyDcS/ZuakocmIjgiP4YDZ3LJOGl5IdbSka1mkrb8q/W95a3
FTU56jyTCA1rFrUFHhElfCUwy83Wz/d4/rX3u9tjF3SNY6ysmUPPLlNA4gN7twR82lEZ59oWr+vx
nre90dNIrK2eTUJe5PrhLhQM5WXPLUdH6WVJwVzT8WV/0UHgJNqWKQE/dgQlcMpqGeOImZX52ZxB
d4hxyvrvYR3NYfKUbMQBRFYoEBRKBU3nrWSOxp1dagKT7QjnVpVga316ql248yiT7s09NzMhtDBX
OykKHP3wpVXgbLL7xfBibR3qLe46f2W1gr7Ki76iV08mazUa9A9b22ZUoXNJHr4dtq3M12ZadpJJ
SKvfOCg5QDr1A9Ylxy/76obYV9VgyWQMoHt2EMvQ1U4AZAyvLIq0LaUxEHuKLrKzOdcYB5c+JZxX
LtkYSwsyAuRjxFwGKzWlXyrcjTm8Md25DlI/ierQkeZvCdtIWCJwYPSYSlXy5vOrG849RkEvceOj
6DARN61WbPSfKNJdZWDLkp2L4w6hBtgSM3/vb3hpfeGQKEhUOOWrTwaYWSAk5bpPTZgme7CpXx14
pVL9zMTmlA7/jxrkGkRQ7pNgYt6n051J1XoJuJvdj+m+LyBfVapy2effYfIkH8PkThumN7bR8XCb
ALy9uD87Ve1YAtc3LdO3uLSi4wuv7FdwURgO5g0rB5sTeB/J3ZgRPWoVVqVQ+9Jey2liDpqAzm5j
MCb8q1JXtYYXnogMzD0FOZhE8L31kDg+7CRtiDFR6AadNUwWtRzYQPO12Mni57jzg99JEbM4LKOE
ijO7WHeYi7BNndDfMW29kZVWGTuZ8ZSCGKvsUcJLlOV5M9+DKDgVn0psHMV8xiHnImBvK9AEt9NE
kmFYQ5RCbWINtLEyBOUVWRNObNtzdd/0ocosZat6nWHwEjMuzz0CKVa7b4XQpS/Si3z8OLJdVSaZ
OH1tTcSL51rUJ9SkcXhYyR33q+CBztqnV70xr2X12Uz7WeVbyds0y/GDDoJEBdc2dc+goUB+VWT4
hU5QyoglUyWI1YSh7VljNUJ7XZNBCIBtU46BM0CHHP4b5JSUfAt65grS50kxxGm/jnaONeuTHBcv
HRLuUAjlGslSXBT01TwAS+GJeahdT4mOHxa+MLsPSrVlIUsmuvw2eWvT54KWuOGF+C2xMlryitlx
wcoPG74mOuRoE5C3piPrEEl3L7LJbtawQOBJTUkOCTzy+zWMBcePJCm6DdW42CCLPQCLRH+OYRqZ
m5ItlXGzN7lBMnp/ZcWRs+PxHG/Fo/2+HepavjAgN+Is4+I5ROF16mcDQcDbWF3lcg/AKEBns3lb
/ygFwkLG/cjHLydfk6Xs4ztcoXyvYqlekB8IF84S9yzrTWAX3at9fQYp53xpo02glBG/9MADzsdi
echWeEI/AY9LMuzcEqoyssM5uZu59AkxeQ9WecXLLNqbLgJJVyIrMKqSMhLbcCwtQd+0yp5zxY4k
t/FrnOzAZ/wPRMNKCd+4SkEnPYwpnb0sY6iknL+qaT+YnqyJRxJm1sqY4t/1xc9fWyF0En8hasZk
z1bTAR9nGt7E6TA4keriDbGUrN7yP4EYxOkp3L/V5Zl+7nYrvXtTqpt2JMhcsC6ta2im/RU5A2BJ
6Ru5EWC5KT9AWEo5bTSovOLuL+5F8PuiQrNJVpy5V1or8GrVHgR0smc5EtOF+5A1yFe9wrC/C78b
uq2NLA7y/h4m6TsqXZBodxyX+jCd7kRIXBy1NynXylOBqNyX9fgpjOZBE+8BkuAyDKFFmQOuxIdf
OQ7rfzqbj5MiHlnLRDddrTy82aGLen2Dk94ZQ46LppkE9gYBaYF4kn1/4F2vvUTBA2WqVTK6zv1H
J82VvaAhoRHz4zQ6uNqHGi8oMn6ycehZDdhXPKBkM2GEXJO+eog4BYEQrvDQg1vuZ0cC2QcwrSgf
X9rTncUuboU7FHyqmzEeme8lsRj5rUerCJdAR6RjsSF1UAH6Oq72eriBNkFvWOOxJqvZ3Kh+Mchh
9JwwaWbK1Zq2P6IddGA5Bc30mp1GDrbG3Zce12RZwNtvCdhBANe06uR2ZK1Ol/n6KNdzTC4LUAE+
mBA4YCb7cJyGBrz8ZSHiaI5/8IbhHKX/TGyyQRInUtihHWwJHGyEJOwc+Lr2BLtRcPZZLBwzQD67
ttNENLEHprl75WNQKhFXs9T5QrJ3z1jLSBlidnENwY0Dxez2qpBCnKhrKbj/C4PxcGDascZEDu9P
hqYbTCXhAWR7/fhIyHTc4ueRQhvuEnK9DIMUCXY9vmnoJ7u1c24m2Ab5djzU+zmNA6aYOU9O9MmV
wdmPE5M0h2O/6/70a9gOwsvvCAstqAnudpRiVKMwF8O1bUBbrhpMf3q8PbHixRUCYI97nikssdq9
Cdt0887tdXOfKWddHTjrHQIXeVH3RTuxtUqIK7NRSeon86/G6YQcJcapJcPJzSpQQ9n2AzQckzPV
G3LbTbVM7XVyu65Xg/tXHeFoq8FEFlOQiVRnDhTNaMDXNb+SJgPlNmLaYN1ivUWGQujUK2UzBsYX
t8myBz+OheSLeOBPlD33vpmKLVxaqdLDc8da2v/WlfmcjICkGfYGPbZLEzWZU5Eelp1zEClbZd1a
uRdHsF/hCUbb9R04W8PMNuvQwAJ6+728sVwcxSMwCDzbQShqhTsjtEi4xW6sRBlwLQQZKG5zd05v
8GfNvPt5jQ9WFLKOWBbyn9THzFv752z6wHfTK9x3P+c362/etekaycpYY5e6zCxqGra9M2zOqaFv
G3wwO6IQcu86O/l0uRdd9funfqVUH7vCElJlxB2tdCb3ybYtDo+imd58p2uRPxCDBrD0kMMRwop9
mkWzLFgm2Y4odDKvaiWdVfhpJlI0g6Al3HijFDNGerEwORqE26Nq63Q07gl5odmbGUStXBhv7cLO
dqFBBnlHqDjYiaMF68v1qAHibUMIkfqw7/JII4K2B+3YlkAHOTYsnqqZod5Ef0mvJAcUvWoWEUYk
llOUzg75RipQ+EKje8GZUbTg7HRE89/+Z5HI0E0EbpQhPnwVXpbNr2Xo72mcj0+prAwnlSfMJmjR
MxMcAPpbzzH0n23xQKKowzqpDhv3S6yIIi5OSk8J0vjrQnyqbLadpTEO5LKhTk8kI7/NGfaQHBnK
jVdMD8U1dyjBEAr7vIovmH0l3Gf3l8QFRVL8yPnO23Vx3isBNSNJgaVStlG/UzHQX9XbvcZ1Xjkn
XO9PJgfsMtF5yPOu8Z7PNFXW3VpbBsixdX/9K8WFalZpnA8dWDtZgUSGAScjHpE5Ij0OFQeZSLSG
rxE3GK7c2mddyasIrm9fD3dT6EAoHOcGu7Lx4KA6bdlSrD+GmBJdPxOeHCwyIk/x65kx9Ioa0w0D
/YwUqUAU74irRcrCe5DEE58zsszMkUwfirjuTKw9bOpWKvPkn9yhWYonXiOEdBDMWzMh7fbUq6hP
+GVYU/ZAIniV6tQT3pNZViYYVgnsPq2vxfgYGv/wgLTvP1w5FmNfoHFw+q+qQjm5fg7EfZCwNuMU
N160Yv1HhoPUJuXN4TI1oim1vfVNP7/RS+l3HsZ8FNkgVFrcfaDHdkysvcjWdOA3jwGzQD6VDxZD
evGT1yQQJOOP/l+sExduY0B0+xQzi3uv1hJ3hJ70Watl3viaE1t9tQm0lSeTd8GPVwuyBKT34Qj2
7hXBs26p+QjIwM6YzxysLz3Ypdhps/i2SrNY5gIorMb54+3vPZxcv3VGbWCfQc3UwOevtYPYiAQW
f+At1UUXWiMl1yrAMicrbncOy3TeNG+pWEdblv8ZDi4mAcLBtswxvx59NCfW689oXwee/sZOyMNv
lIEh1HdJWc1uDQWb0bGpKm89aUbf96OdRYv78gufHqQ6SYP1/DgdTJQhxl81smX3aEcHHdr3UoI5
E45LeVgJmXStV4py9K7x4MD2Yml5953OA89jji9VLfP7JFBFTBoskf6rKfTTvrN764vQJII6QDVy
AW4wczM+5AW/KWuBDygkxqxQ1+t0tUgOSy1esTW3PwJvL2G4aBGIYNEqAWmj+2IsoQFWGvaIk7L0
fxUnK3NEeGIIYYrgrVDu45355h7NWwy4pjPLUwUe+tm4msfswaO+pqzF6Ns/fOWPK+6BAhYHcWz3
yOWi1fJSEpf5khIA4PSE4I+ggAYkoLysOnF3EpRVlzp0VC/NuFk8/HVI9fceRnPLhDpeU7P50SX7
Y8RtcbOoQl+C3ibVHrOzeha2m6NHE56Jp7kWTrZY71sE6laxqNMnEr5WVa1xd7+nSDP7nOEO/one
YwxMffx2uvheMc2YBepUMS/lougUz21v0S07sPmlr1MuLbY+jibVj944ZqYVdnrPnN5Wv9IeLXJG
UxUpQgQ9AcLBigH9zUNu4uf458yULiIbboe13lSaSGoLF0f6nFyv9mJx8kkBT6egWpz8oDQAA7uu
03+MdUHeiUn4iYjNcRDtr4NQhm5S33tGs2C5mO1smDWikTnZxWTLM6jlha9uIgVWsEA2VAlvsj9t
tb12mkIiT8QJw8SF2SQobJSr4BbJE6oI/9lk3xBqhHVyRi+KWb99OAsZUGXjJmj/6KUBLX8ks9BI
QQnmfqA/4cLmGZoMETg7Gd4Udg3zWTDnX7eX7HmQcIdLbzpL+c4KBGHDjlloeDjIDdLdkrBk1hPc
c5WLRDrZd8zxwE7hJoxPolBQyOQBAPe4ApA9RcebvGaJU7zBO8lt3XoMGNiEmoaagcpMyIbhj07D
PW8THl+Mc+QRjMYr0qDY5oFnn9Cqzc5OwXBvmvUbRxfGSifEGh10r/ptr/BEXu+dFvAwOWcQWaPG
X3BQo5R7MOv4DtEl5TF11UQRvvFKqH7sN1k4jJrYhnAKPpoeXnu9sAYuM/FRc0GPXAW/qbthmVHF
90CDMdKpuLOzzqnTj2c/mBf5pO/vnjEbHHZV0msX7G9ggWb0CUtHjM4s/uRKLPF3PV7WyLl8qTmc
JYJhVLKTdOtGNb7PBVwKQ5kbsx/0EIbLsSop5OXrb/QCRTmgzHG3reIMcFVzubMlXPbnx2hnjvjk
QjzU7fixb/nO9P++K0FpbrQ5dZ4DhFSxES/gM2yhnHGpBmtS3BRPyu/v+pboLqytWCMJx6msnfAq
0LL9KAJDtCRsvh9o0z84Lcka1XosRgqwRVMmRHcndT2v6OdkG6xNsLQxctkhQS3SpA7Xe9ch13i0
uYxksKSmJxlKj0rjemwW0Uw8A2ec7nIpHipnfH/vp0V2v1YP/3bMHBJY0STjvZteYpYxUiqF09Ua
g50RQRHzVJIoPAd16yyENRAx/p/FSgvTVl3tLdjcmUCePgV2vmzFy/ixxDVtKJwwVPasRbNj7dEb
epXvOgLu9Irjr9KOj+o9RL7dR3v5d+PnJ3ndz5N9XW0EXzXsq2k8Mj7LMCuPNWiiyaHURqyOPgZ4
3Ft8M+sXN/E2sOhgnONBvKLttRYfN0D48rIKjqogWsbFN2Mj0PFQ5Lz+4p5Y3eDXQAnWFjzUKsqX
yaZR/RwqT48LT9qVx8CATYCktYJUnfXPGuVHj8fNC+Mok4ZYZBfQLTJs2dzuMqO7HI+QfH+F5Y7p
t/0koabzFifayGZ2Z36wxrrPyiIFVWrmg4DHUAKpnJbMf2wyqzGvUnRGb4p2+PvSx4EggsJnGlLp
hoYj7orGe3rXWGjgML35kPzJQMkDzJ27wJJU5vPylXrbwhFC49KXeb1ec1BaQIdMtWSVKOBELyEN
Xg7dhf2pehv/Qoq/S0p/ip+OZm/ubxqSfRajMJCm8B9AqtIC6V6jhmj726fAkQcAgvARmM8r/mSN
gDKuRZ38kaLuf6AA4vQRKxdYfCWy4lCWbPG0H1xab7ZHivo7lG8Sx5rr6pBOE7FMcQrvzyVwnKLY
rJtBN0EV1iFMjvQikaZ+fM6mOpG/0hCNTNCtIJOZNcqsNrcFUjfZsPQzCnlJEGpf7b1o4PsLG0px
/wYmwRDuQqq2ptJsSKKh0ldvGm5fammuOqogwSAW8/0kttMt0lXvhDUVEcS/Eom22GPQfSci7FeR
j7vvUsn5jVN828bi5VdSdn/JtIoZf/rxY3SyCVS9MbDB88yCX5FwkiRQeM9zstl5fIIHmvFF/G2U
bzzc6sgsgJNbnnPfBKPmRJ4a65ASSny48XOSjU1ra8niEHmqgRCfPJSjz2hJtZjQu6fUwYQpvLFm
m+k1YhKq+186YhFyNASmuZUOvJLRcKlskYgoIHtY0yhLmScV0FW5esROoIr9y4kjEY/aNItTnN0z
5gDGKuSVdUx1sKWEtVyAYA+4qdXqRTypTrfxoAnkmKger9z+OAQ6kFvXYAxIj7Hwff7JSVw2XISq
7itRxx+pOp7gKi6+j+YAMh7ncNeAPu6oNL6rFAcYtpjncZrd5JsxaettnJHc0F6G+UkijmTxkTqx
UXjokMBsBJF9v/jKSTOGMw+m8bssEN4tLiyR68UPt25WayiQDScpQkzHAcVWbRkcZghJ+DfOxo3h
SALC2i3D3rGRYPMp1VY171AL61dOJyJneHEZpj+iWXe2JwvLsG2QsXlred8UrKxUyqgoaZuJw5Qe
pWojjmSftExF7sqsnx4vYB2iCGPVZ8322vPtwulZQ4/HAl+ESy93uAHw+Yd5Dxi6KQzT0kNQI6qk
ImrG+GyCEbww6YUWvDmkEaPM/xIejdPOY19KhM2Vl6+gscYU2qFpOAW55RyRQE4o+kWhTpD/hfme
RTkLfvLZknIUBWJqrb/4gTcTkervYwIxslee5zYmlH7DujsBd+B+ePYRLdqHaFJ0VYYxl29QwQra
pLQbYFd1o7GubB4EOPHtHyt6hFfy0vKpXZBt2rgmp/NUzhymE4Wq9I2oD3gjtJYdonUl7WmMPoqz
IVyxNnLZPuDfFlfgXbzS4inqfN99IFfebUwZBE3wqwnqQwh31KCQeytwQkdl0SThwL9EHjhi3pAV
gYAwDwx6GH5FcejhVr9CqufYfqCi7TX1RkdnsmDbcxKARaeRVQW+sZLVp7OnQ0Q8/FZBnlgl8+tW
MZ/F+crLvnZ/wE61doaWopNkBcojtEKlVXphI6uTVrjkRFQcoLQkpKW8ir+cLFKK8B90Ib9w+hZJ
Zcr3Bb2CpU4ZKgCB62oArku+ejJooexstoy4aB1klh07FEwlQYIBkSn1sXGxZEtASuQ2YBSXQlxC
KJr03uX1sN9qoRDOD5qZ6XTm/bQzMcyu9FwgzXZc4bZWxnMl65f1MYRTqiUJFsXG/FgJ/NTxUgZV
Y2bV+boZbUR5aaJUJcW478NbMsDVvB/HbQSSoHqX2AKFt//erbZmayGKP+w4D9KoSv0q46vgfW6I
ITyq0a8ISZOhYenu9L2XurQpd42dnG4eKHrNDJzNHr7uQlQqMJCDpUKL/d3+GUj8x6E8l0gib4Yx
NS4qRyD2fUNb0fIwu1zGmIQtFjkknB0pj9TZw3Nl5poN0hOvKrxRbphI34778IvwMIMeHSG+N+Yb
o4TlhMdOsGPNl0SWDpBhddWHoPEl9jBJTfg8RWN24vX+QcXEwQHIrxV0P4q3KDAr7x96tJEnzL0v
2rZ7Od3klZ1bywLeDOWOg2Byn6TNsUeactu5oeHyz84F2tKa9znf6jbaFQN0FMMLEqsLsgtE9XdE
Y76iUNKLZc6e7WGrg4zGOMJCzLk1GZ+lAo6XICPAg8CdGTR0kMVFgfQOcYvwjsDTIskfaRJ0wy8u
L7AruJ48SunUWO900gbX4e1dSn4qjb5caglr1q4zvuoRplxOHRC69twLluzh2y1+tBs4u8n2pZBI
1/TO+x5k8BQKYMbgEVT3/xEqscn1LR1blw7OKgdndsRmYFDMkrQOE54OLTFRxtbki43P1Yo0uSZV
llkuQXdQ1kWVW4KP/FUk7ZH8N1uKuQU1xPJwbuuC3RehRYASNC4Ru1O7V91r4DC0pycsy79+LaOY
rXpacLSNMHS9VRz95EwrF5erxmQbb4y2sjFMBgI9EJy72L3LepaYpk++QvImERELPVv6emycOJKf
C4FJPakO+dDlHdUeW/zIDY4JcBylm28cC/DiCt/6y3Pt+bVc/vZRiaN98blFZlBmI9V7Fshtux/q
SdatXIaRU5xWbZyOo0ui+HjSWQxdDTsPr9Q/pMHV6M4dv6RciCHNxP5z2MkU1Z9xOndWFyUhBy+h
2fv+yBbal7JbAnLajJCvDlfoY3ByU49klprahvf5eZYIbGNbQAgUzIYGx7KwrnNbovTFatFFrNMe
Z5Mt4h5qPB//GiChs1rKOXqHB3VcU0Gu9rRptjn+4aohKBUIBP9Fu8pP/Rq338PfH8YoxAHoHThI
s03rBPBPiREm4F4FGRVz3TLJbYczvLbr9Tbt6Z3kq38EqzNl8T0jVO/Sxt+ySdMNiGgS20Xl0fMb
OgKglFtB75byW7a55NBfMeZ+AEN86AvHEcE8BE40nfR8r/KfIxPWzez42MtLaaawfr/z3ajkPW/D
nl4k0vlKiDFl+Wn8lYXObyYgHmtX8HzKWyPCgVFBViySRXy8NAA1IMvedkdoeVwVehfXyHOhMxkc
14iTV1bRj7yxrsAiBd9mItRJofu/ZG4a27LlNJNelKJqItiKtw7ywsP6H4SdlezdfH2WMIDS5DiG
h3jyjjBZApF04WN1RuRPXk/+ynDt1Iwg9OMT2qP2r7L7GUOEXjrQWEeVkmEvCF6iu/gP4v7OT4UF
zAixP5DzYuyA0G3ed6A/pYS4a+f/1cnJXDZ4gwZtVh1Fm1jXLrqBIEVH1keiPMXBKqmlyWFdhcEH
cTrXwOnrmkxlOccp1cfNXTjb+6p1oBLVBW3bRY0eK9R8VL35O9gfZb4nlp5ak4gzsLvZ2zH0iePA
Yl6XYhAc5oZ9vvn2N/a1ggmuHg3li1+xUN58liq15JgjXen0HZvOwBfcCbCvP0F6ZsjxQSeYBvYP
snI3FBKz5mszohAAS1NBN+GObF457woivpEwYxn0e3n7494frd9qizyTe6OfJvlyruNVNsKtAcAU
zDwCIBAznEv/T+u2ECIfFm0bjND/E/l1s8lmuk41dTA59pL6yjeHdFSbRNCtQezPMgTMQZth/sAo
tXMLsBGsZ37c/R37OxZM9myHRLB4/B8W5pJIby08Zf/ZfnVfxPT8wSXnPSwhTp4mUfyWy8zvicgP
k4Oi3uRPd0eAY4dE9T8tvrKK8FxGJJmN0teH6gP54340t1Cd19oHFSFyg1lEZrhqKTLPbQDKklLC
oZAg+gNlv8Z3KR+jFFGgmrtJDKEIMR1gKBt99tMeJ09JFV260dPHIVG5XswGTWPqTGqvVwRfCyrE
IBMX/OgsLq6S3uh9eM9cnOgHRVdHDwzb82Hv7PLJTplfbjIZSxs8fjh3RBN9m/HlYhaxQLdXu1+A
6IJrWow16hh10qgCjunhikwXBsLUuXy3X/3i2J7/i4jPw2i9iUuknVSco9/TTD07clI+MBl97gqa
6KQnSEuE/xRWmnsOol1nv43DjXTH6XeeVKCteCywAyCxy8oGg6AkfjZ+n91Y17TseWu8bt4xlfia
+1JErbqA3OoTCjkTie4s7Be0Lx2/PbgArDy6uLbHr/sd9O7d1CAdFZcoQe45t+6tMOhtfOuqbV7O
aGYtFj/249C/wNXYIZnREH65cjjqIfnfUlbbFQpL8UVczLzwb+STlxplpbtWLu5LaHQtBOUEgZMi
IeEWl7q7OEpV6a0btiNNSbATvEylHMNlyNhMpZv+WykX2KNT2ClcmQryZI3leXqXKJkfDIM9XqKT
QCMczFYiSiTZORcPZuIcTvKq/1cVmSKNQkfmeJUZkROA7sUt/t4hBKBJcB510EsnQxpQZtdTUi2Z
dM0bJ4Byd0QkxitMtLgOLNN/ANsAEbEuFMKeRuX+w1NpkIfFPQ657clX2YPBgfxye4oi0ZiLWjra
23v/TCk0MoJ2JASeEQI1nJGg7fCse56B267yZJVqyt6enp4dvzTLiECOnjLhnTbWNMJRw9Kj6/xj
+Pvjk/O3tlfr7dVbUTPd93DLmou2EECcwhkiggArYO3h/r/uphOfNdgEgQwdMKWZO40eQfLrow6d
yUEihmbQOgiAvK4fw7qz7lsm7/4Jv58QFnvoxHB+TYYu4hYCgZwGsuG8WTI/F06MDdm1Tny20Wyq
E69nU5yvZ6KDeoNoz3ImjydVWM9nM/H/XNh6YWtx/wzGc3WNG0o7vNm3QxPSQVMZChfNDNVqtltW
8z8XH9n36x4Hq3tutqrMs8TONecvvDdpbBfAMuX45Fyry41891t5X69FTYRPilsoGOSnio3IKH8i
3zNkojMEeVYSu0/L8YWHkMkQGG3g6d6S8/kgFxdb7Yp35Y3GuTrDsiEsjUzQBrQ/BMWGZf0axOms
9JaajAE7AnlQMg/7LrrYympirmmG+z5TzmeNwidbf9SzTvfLA21rqmD2rByYhA29rThQPVlQq134
RVRqQfZPzstBppGCRcOt0SahSP9I8J3BzUqSL4Lm9MuCQJKxK3aJ4v63N1cqFTz7GZ/kc31WY9vA
Vf2b30OV/DdG1NOFSFcEUY3zH9ejrHIhJ7ke0l+OOfIgzQf713tho9C8cxt1GHFy9XxRbG1pPl//
i0STXelQmVrbXLvtBilPV/3/jJnNi02/u17dS01nntaTGL3AgBgkf8h8gk1OAM27RDuDJs8avUFt
cLBsng7Gx/YnNClUX8Ci0+EHQYps9uoDWpkguDqvRY6VrOK7rVOZiOp1WroNy6uRDQFrB64u2M+6
xRM23WzgccHGF3Fu0urAxnn6UN4zLV5ddbY3QJsU/98M7tHasvWJIN/hgN8lKQkzLqiK5nUOKFrd
OfsJ1AhsV+j1dOEWneOsoLxiexWaUgX+2VXwAkEbjQNRpWoRAbuFa0jWXgBirT3/11T5QFxkUtkw
354LmXO+9QNGbGzrLUO1nCD1JZSyZzwWiE2qQoXHojqX0N6uHnovo7qsRCrRLTTt1OKFQoLh4AqK
GScWFGJ+wh+xKjuQ+GDvl60bkKbZbnJyvKojF006jMvkrGdTmHnT12/7Q6HXiN/YOURJ3boN6u3n
Z1b+FZeM49YG5lWYVx7MTUxpZM4Lt/itF5ii7F0ZCHkhSzXvIxEAtaWjxZIRoCp+wEbDTlPZi3ek
DW62Qyc4amxYGjFVOCNAgtZ1eAJWWsRrtZcQG08DUMwWCyu2YE5BUADNk3KyGXeWfLcMhA3lqXce
gpWit8/SJJX4dwWtoV2UV9pRl1INYjTlhV4gfSpdVlPWcWKnJxzYfhaZ/FBCys0YrMabwXJwjGln
xZhcNVhma8GAHrD+iAZ8XifdiAMISQRL/nojzRU/yN3Cnoa8/8ERqmngREIAo1/K2dZenbMRi8QJ
ioJwXwhROISNB7JHxNaikSCG8CVscN6kZFxjBZVWx4IqCWBpdZIwFIQ92zfMZqbUbmNZ/MzdwLI7
U9WJsKJvK9Ix1konH17Zwd3l/qUPAL0JK7mi3pTdh7oZT0bSpYNpucSL4BXziVBB+gGO5ft8LkAf
ZLVBIUI6LRKQQuozvZ5rKjWTYxG1prTi7JHwmsX03GfyF7nff8PiN2Xjv5DM53vU/gtZjdDLZ9cB
hcObYKrV15Le4ITtTRzHskgSsCcn/CDt8AwhmUj2uNYqkr0A24VTmaFtokjDaROxDorTse27dZ10
gZ0sYxkjRbusPQ3hvQRWioIQKs61LLsQMmZ13uAn5UssDqperQTS7OyQeRinCoseXiwiaoq0XSHv
QDwdbdjilNgFjmDCAEXuZFI1PVGmnLJP8FoWh4Gt+2jufBmmeiWm8ECu5WiaZzpvf3l+hiHpnGPi
3ZQ28uuaHmVkTGD4eOAI9vJcbeSVPgh1IJV89BArkogz3PopszjJAT6/tPJPbJUa8QVGiqsuJCJB
+V66KnnDO5kyCUWPyvi35koOO5pDcl6s4bfFxOU2U32LtIKVmczZNhuEs0uakJ2o6wExirrUR4Xf
kJZQXE7Vy/H+yQ9S2YCV/68xK7ks1V5PbgZHLrDjJ8jcl0F5XXaZmZ+HdWgr7inG5AArRAsTXyyY
rPOea+XLw+LVkBPJDuMX5eC4KYS42cSSa9CIVYnb3SvXqZuAFu2GZsKu1W9rZ/6i8tlpXduQndC1
HTXE/KqAITOKPx1sjwgXjpbtkkA+wixWLJG2C/6YZ6LpUALEu6B360WK1ka+zu6RIatExhQ4A5gT
965rWZOFzc9YgXtz7pnSY+UsV2FBD8QyZvkTWj/jsGKDgFXKi/j9qHECNX29Gb2ukzxSBdRr350l
pgQ5BLLy2LJwn43PsG2RIRw4dBD4/bJfMnU7PnncK4trw3TTeR5hyRxwAVPCNlcnZyaGtj0cuY8c
SG0yRfaPWXXZAdxQ5CjqA66epHu+VQqk1Ie1SKLA29Ogxmd37beGtlQX/e3IeXq/PZVzcbMh3Uw/
t06Ga26SgC5n2nCUMOIeeR46PfxV7ChgVYcCz9bW6LbKjIBkvUeZGppzwqRPojPshmGm3WdXe4z+
x92XxeCY9iw3KRVVMmPomxVvJ4fOLCQWisNwWaxtkxCuRIg8T4SDD+ogNuaAChBd1I8aWJyUoosm
Fj8NTcjOX2soj8CPeQMOdPh6b4uvob3Snj5URsh/rwb01gBMy9nGDl8r1rGIgGl88giTnjepp19P
9hDrAqm5vp324qdI7oDpQnDqGQM72R0aLCDs5PcS7geS4Zxv/4sT2BJcp/icrNNAD3FLKx/LDO55
L8M92ksm5997SNCot2F+Amp4ZRAZIt90g0lORt2dhjm+U1B19rNJa6gTHVBqD54gIBS2eIIjxpK2
LJ7dFKShqHHblXLR2LF7S2umgzYjgL90EXEQynntXwiOSLrTcTKmUZAGFBlt1PSNWlwM+xYo8DCA
dUsdvLS87QVIIBLWRMPsyhn3eN0f86HSZrpY9YNW5f1C9fQymazfLRwigTGtg9k98vK9pEMN0Wv1
gHMuqjvAtiUKaY1MozkfqG/Eu5+QrIAOSIy3QcWlQ3u8W+TCOvQtbyZKCrxEqpVbZA0eieuL5mRu
jgGGC2B2AKtf3wP8s58FSWDGk0u0Lkxl49msKasisUOox3o58RUXqOnPGu6bjSYWEFRS+qb+OooY
dX/7hfP8vkZFB+rYVgPNIbKWumcyNJyE5q0IKt1ockm6W5IiaoL4UOwRd48Mag6T
`pragma protect end_protected
