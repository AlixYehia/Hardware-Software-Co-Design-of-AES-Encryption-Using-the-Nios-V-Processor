`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eJ7WPHKo0/2FHQ/Qp9gBbUNIhaA3s8hBFM11JCUSyurGTR62PVkpsc0Rqrc0uuWf
VLceh7O8NafC63cMe6Ba/lnUJvWvGH/4RXqTde4E+0pVobctRl6NYS0XCePNei09
vetJGDlcMTSZ1uk0Xg7wHwQyxvvqTeYrmjQYvuU00yw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6640)
RhP4dAXtnsOGpMp2vQhJ2/BrqrOyzP+6Wd0l0Xnmkp2mUlz1iGzKEyuWVJG1AH0C
/IIcOwIBcNmIe5EaKqe6wfBR93B1KagPyohMxfcMHSY31HWDW48JNBcpQWwJsfEO
oE5TVwY/JgHzTpQegxyWd3h96JCQoUYz1RLTnCl1rRWLOJc4m8rn4VytLfuLkDCp
F0TSIUR+eAqgeSHsdXkZ13+X3lN2hz2JxTEgojesYpIrRMq0jkOogoyj1y/AU62E
5L1FJB/OuUFB7uZJgoFXDQ12Z2pcP5CLrydRbLMRBkPClg0pk7XA19S9RXfyTTk7
Ca00vnBKgOfouVfqhGbHNBIqN+hkhCzb7GN33vMhrtXmebvr+CjkicTY4jEMEmG0
by5dCh7Rqt/QogMo7/mN2k6laXudIrEVDhFXg02AA+qYR2OVqLA/VmGybT5hoK9N
SCk10bpNExStdJ5Gel8o5bNPskGboqKzW5hAAjn494TS20FGjIquDfu5CYXXT77f
t3lRPQFyJBEADyaM1eJ2Hm6WLqEFfoOcZSYDwyX7txJUGVf0sfKCfhX4yuXDApJg
0OV4Z5aLk1ZpwahXRZpriWY1d8mgJM1RPoJNNFEc6yRAcTX7KdRyRVwCsOhPkRP3
ULXqXx2Y3ArbJUW1uOPe0OeD4BXEWWqC5CbbzonX2JaVy7uHDA/z5fbL0RwfWJva
lB9DkBnSsD5LTzl4PNQ38sAfZPt8SBzZHh4dih5iOoKd5y6l+jDfxsxe+DXyaGVU
WwxcbGr+tdrxkdl94dPX9R7RKqwjnZO9sbG9ogZKTnh8M3RUuzenjmmmY07QcES6
pljhjfMelrKmmPwJgXllXIZAOuyldAUX8RK6j8Fu6nCGFi9rcOPEyZpRywn0kXkI
LU6mSmVMawMHW92rtzaKpFYmn7XnARdEjxq6fSlEgxFmKhYnOT/8wUYkjwBGmA1P
EDwvyY2F2XciHm3EQnAdef7s7VQNr4yco5qXSrRv8sqfm8t3QUPVTYcL+0b6KNV9
p5AOff9y1kgoMaFgpVCyoe0/WagJ2DKK/mbIIG6YNusVeVzLgjYiMkTe/JQqFSTb
9tNmJUhrfv3k2vuBzo4D0NJ5ACo6fJIQmz75ald0ho4LF+5O3BqKLUg2F+oes6xd
iQTYdXx5o7EVjCFpj5qmMc7axCBpPQfg7+vT5j6d9IM9t5EsU+Umv2ffqBVlxFQ7
7VYn/gFSuwl/m+Hc7scf8Z83GppcXvrb6SGy+XkgAW+YofDlYHD82Ni70VHTpk0F
Qh8+CDB76IgpQrJhoVqI1igHUfOq0cZgkWMQhZ16Bbd/pgSlcEIAc5HdKn7i6Ggr
DyJyK8P9mcvZysYYLp69m4VIhTQhJsVJTkco/YARUU2yvy0AA8SsVoE09cL+gYmJ
DJ5+7w1z6WlC7+Xtpqwt2aeZprVwaY9zT4hUN8dkR6Zx82K0xE5TFUVENyyUwUKr
sEXPkv8CeA6Y9hGNHP4y6hrM4LZfXI2vlN0uaRbaUxRH3IUJe416MzmmgxHkbUNA
T8/LAjkuuIADpLX6WMjr1LSpm3wezhIE5mh+5HMfDyEud3RR7KLABmbwLeaQzxK9
Hpc1Ftnkr/QjuQpP9xkqTjUSukh/fjsWqC/h7sq3Rye6Pbx7Lbcpvo3eaBwLAbqC
IWlfpsfz9bZzhtUww7/A8n26UzJrJz5iNP59hnCOsRA/q7fMeORPxT+Gea70GXb4
7pQmQ+zDhWmKPZz/pPhvLDj4p/+JChJoGzevESxVh9XeawPzaYKulDcuCF7MKTEr
BM9njNYotW7d+2ThctDebwu2Gn3r9Li3QvZaP1ZlNs5dvzMnRhWTkJs84s3fUSP5
2zs+rVFfsueve6353QRNgJIQFKcWqt7okSEXq6ilFv9COdGP+PTfmZ8heaTHtUWn
/hERhe434JVgtwPsTgzLPvHLvouXLXfPBNvRc2tjpaftXGyAfWkVxst4u28zSvB4
lb3gvpzhLo0aleFwaT/NkLE5xhq32XWvQmqLU1hYZw/ro20tsRtHnqGrhF79Dsfn
ymV1Lb7Ldoz3TwpJq4h1TJXVnX5XwLU9D9vjNNcCMu78N2XINZKrphaAVZr6yN3c
xbdsUlZUHreq17ykh6sByTYwut03NWAcLDqq092JDOiiIUQrOYgfK9F7GQ1G+FeZ
g+r6QtWaDMXHjjGPY3wZ4SOjF3ddQVQmnpvTtsUUfFfuc6fQqu7WYIoMrYnCEFpW
P+T0iZyUs5yfeZpb5xzMNFnXaw5YTYBXedDRVOU0AY4udwIFSPmOjvT90zmbT7XN
D1m06iM+ElfihbugfmvlltZpPAvmRtc9AgZykRMG7ILCCsNARiZNEa6dMDq1e/p/
FvC54pu089enY8GgbmlfcVNPyor2hy0mKFQKduAO05J/Twg7OTpov1mmliLwxkWG
NKEb0CT1suU0AwMiKa66axPkYwxCNU90TLL6VAAu50/TP+6JFACpCZrztdYxXXwh
6fnr/TTcioFwlq3kJgIj6wIjCyuh44zFNXQkwEU0GIrumnYx0OLVQL2T/2vNPXWj
Wd1jHnPHua4HvD8v0vBWMIVL1jtpN9HOocTbpfByEB07u5Wg0AP3NeQZljIvO6pU
Pr9U9QV+xdwOVHmuwCAdhxQ+KPPTHaslAVdvd02LfYO3ohtIipxHrg+36rN6S7Vg
oDvWG5dEuzIJ0fij04zD7+AtDB+KS8/3QmwTXszNFhVCFHj+lKFBJBnO+IDqJHhN
tKwUpFdRSNc+xNVV/WRlqgMWvQKXFo9m3i1eoZrZenf4w9bRDluwRdiirPmhPHvv
lqRzMWi08AbxDIgLWjVLrI1W5h6B/O0E5DmuMm2mh/FiBDjZVLofWSMSWOn0Fe7Y
SvA0w3+KpK1SpEWVFhuOewcOcA7HWOWBvPsZ5XhXIBtQfpfViIOiMlw8Nql20Jns
arkYf358s/9erKjqlk5T093GXGA9XPNF3Z7lcrF5md9EU66ECVB/bw83CIhCk5l8
P2oa7mJzAttHx+eShrR/Y+pkptlvK4Ixdh4kqH2tbbLIrZJfhVqifGZPpnUqH9nR
fjvRCUDH54zRNnaXpBk/HPGUz1FKZEwagH0m1tcepPevCZTkEhqztKSuie3KI2Q2
8FxlRfXglnlk4P8OifurqDAi3tcVqYJqwAvWkD+BNBhrzckxURSBJalX9TXHDzmX
RhN5F+RnEN0kJ69rssKhQuFSdFhbVdLvnEVdnutf8G1vPuvt2Uxw3zs5lQB6Uckw
GVm8g6WHg2iwg9osj8elkl4l1Nwc+Q7cdBTsDBehJ6JRkWMRuSRbK5AOo04U8vok
ziAvN5Kqv/tqo8o8cqBwNpE+khInz0rHkQMZBhM/+d+Ft5UsTgM0b/N9W8+6x5v+
u21eLvfkBB5RiCkccZhTIjmMGkGfR46w7Qdezr5LIzZp+nSTo5pmMyHdu/sWDhCh
ZIB0CmkuanWv0l2mKj4tT8O5YBes6bIo5AG1Hjfi7fbpllXZN1i9xfAf0S/PrhaT
bZGcVpk8Y3+8rI5S1IQfiG4zj1etsA/G6p+xgu9yH3kW91YGWosr0ZP11ddkyRBz
yFYUsHGGxMriPX1s1J/UC7ecxp5IjQFlOws9J2W1v5XQtIEkxf2qaf7EpLE//qgM
IgwMfJi6SRSz3z+WcPrI3KGca1iJZ2WY0xwpKyls5rWseHFACWcDe53gN79m9xHD
4eTb5/DQY/4XYKUIsP4cgu8chsUxXPUviHPaO8jgfFFOlNjDsapyVpB8g3JJgM5m
PWjNsIMvtyQPrWNiDu3yzByxmMF1wfSm+ndLOTe5qQCmW3BiYVLTb9/xiauTYEu0
sm/PBtqC6mkUQWTX8Y2KdxuS1poW29a6ex4G1+ePIuhjgKanGQDXbmVDQDTi/iYv
BIoeo9sT1JXbGSaJP+MApyUKyEGvCAU03uJUgRjFwHQx2muTna/fk9c/6Qcbg+2p
nX/l9pAwi17fZfNoV9sx51ygPMmte5iydNyEEMI3H2aPptS2UsYif4QFGqnM/k0L
Rd+C7uEdWOUzLqLt9Yzj3wvR7nfyRfLyf8zYGsNxBFbCgyh/PObFUVp6u7xRYP1Z
FKFZJcYRPLk4uhMw6QgcLaJBDQ/uf6Bra8F7FII23KdsuMthQX/cfslqhqLqfFAY
0zB35vVsyvr2f8G8XS+XmOECn5Oz0b8JpAi62mb73GgHHXFC3RUME7Io5w6PEe07
5yHw11pAS5kXpz0csdcJ+rTcBmX6exBdBUnkzFkX9MU3u3upz8GwWLpGGLpQdKZW
Thj4/O3gI5grHoiE0ffg4OaS+OvN/volt6i/NyvfwOxzWcRf6gpALOJMlpsFQ+PM
Wgp5WUzgKyA5aokll4dWNbqVnlTxDUMhqF2Jbl7NAIZnd/kVx5kELIuaN3ISYSZn
okaL5H/rQXfjXzxfCYHc87CVI2yvSP6EMLE17BKebUXjI7zzpQY+MoDyD3f4UeEL
3gYNNUAB1u8ozFvpeB/sZ0E5CBFq0oEczo/s3YffPhcHPCeVrUcU6Wo6hVrdKPgZ
Mme0Wuzy1A2ZFW/UqqsQoLhywohs8xgmSBwbdgFENzgQjRwxFrw3Oup7LHyoScDe
tmY9/529rG9wX00MrTDvTY6REjFfep3cLCo5FowPw5DfTF1JCgPvxov3nqADlpTy
KUehxvxe5iHflft55PXmmInDThjOBcJTFMduf8OoY2BIDj8/Iz2/MetjfsjysOPx
R28oTfdvdJbjnZjOcdy4idOphz3ZxjyW/5BbrCEmBwY3RblwD6ITaE1BxodvphzQ
D6sRC5s3uhp9zhm16N35Nvu8GqEybm+aTNBqkVKgnpesXqD6TydZNEkp+ExAXmif
eGrLuwOYWCHxMV6zq+Pdtmu0rxYxpBZTr2Sw3R9UYyr719oQb/3es35SMqiFhWlh
UPp1HQNgeuv0UnPzNrp865W5pETNG9bCzh3QUaPxPQPWSetRFvl5o4IWYjYMyry5
F5mP6uSRVRx30ze1I7VPh2NUBxunE23xfP3j5nwZP7LyrzHEXCeKI3XN8t4LD9rK
gZkQczQqdV7uY8+eWAvhL2NKkM/D2kXuRyF0tlZzRpCPSt/5c6iQahA7DKUqNu/i
oNXrhInI2/TY4ekLptTc4cIRggrqK+w0GosNNuC+emONsW5BGV8PkmsqgN+36RQE
UNpqHV8Y/HKaodqU72+WXr2f9vAgmh+y217N2q8iqqRbsVtBXldZwEA42f6klwSS
D5/7AM8YWSXU/2Z9Vw6dNRhBPyf5ChB3wvZZGJaSsIyw5h9omEBOSloCgpTgrLIR
fk9sfOycDRcY+L8ppvJUjtmZU37G4enuQQQ0ldVJZNjer3W3c4h5V+a7cI1K54v6
uFrItVJLTz9GKP7LTn1I6K4bpQYs8TZjM4VxtUrF3L9H5PCjhx5QVG9HLq2ggNBk
tt1LhbenqW+MO7LC9Q04RuyVq3SW7y9Nd2AqMrjd3Se7Hc76wRatrL7f3zgYfS0d
4k4cpkl7ZworDjKV2ZJckuztNOFoMidS6/oe5iCfJYQn0vdseV9LVyP3wLx6gTmw
WxlihISTsAq6zi/rQ0Y13YG9cQOHAAxrKorQWWZ4V2Vrxk/GruSg/DbXeQDdzwFu
NaQ2iBk7RqkNik4Hp62qNJLhPJ4hleWRtdc6QrFgoTsDWyLn4p608qD+Zu5Ptodw
rMv8sWJwhCwMCT4mqoLM8z4L5c6vTHZFPPrYVViZWz102T8mw3dAOE+6fH9ctLRn
XkBLFEfkIRxqV8+wM/zxh7u9ryqrgrjd6Ex4utVfB7VWMdKLj2xYwy9qjq80mXtA
RNTDHjlyMSfhjzb8nAUAjFEqi40ZVJuouIw8f5O46JmJh006rawZ2dZ8k/mA1+1X
n4AvI5X7XpI5cgQL7580m0p/e9wiT9r3DLTVFtrTCcuEgcBnl2Ts5QL5yNccO5DI
AnSgSypVeOfqEi1NvZ5LpXBpr8WnfKPW+Gy0/0jkG0ebDKiRbuFUx6DdMmqNoe7I
kbesWwybQgcuBSdPWJVTEGgfk2jAw5YUCS++amJwkUaOUF2O0k2Itu1mJ9yzllS5
lNO87hAHQlVFKFgiRNAvJjCR/YfD2ClGxXYA7d3lnmB6hFqePRHZ+YC9WZEWrYZz
J581Ux0jkh78g/xtL5YM6wQUDy/iQWdbsJmPWsYeKngafg54aKKBwzu4NdWMH1sD
LSOBMWt6WhTRQcD3u1lG5FwG3DXKxS3uu3KjGbAPPBpGM8wnFvrStJU9942ktwLO
pFmdrUpR4dFmxvPI62w4KoY19/fpBAWtDQCXnKliqFfIutZDgvKaw+TP/pL/OYSH
+hPx5i5786DCXyTEDwpultvLF2Gtj0rTBaLE0d+c1FzsA9jRlk8msuWL6eIWREBu
YoRZxK+tyE60WGSijHZ3IVQtI1VtpLN71iUkUwBmmb22+sAwcLlRAJG+mJSRFS+r
PHqUlUbwenw2uatQBU8PUZ+VI7aQbeq9eE/NT0mi7YDAr1XBT+wYFFH1x5ZO+8Ct
p0IaPUrpJdfYIGXO0G6KmByU79/3o449BhTNBNO8PXoB3w8dKc83gIeD+sdoUhI8
xEY1crmYtG5eYCrPM2/hOCOdawvrCGEG3TCVeqN1L64tYLJYtXseItfrlHbhOLUC
LWACrdSLM35ktNBH0K+lcMjk061Gs+AgW4pjZVg6PRaQt0LHBR03/Fi456qBol4g
4ubqLPs1BEVfh/lK1ur9u4LsNU7/dGkeY7CHBt1yiKcOxQgdPiL4tXJSo2sHYmb8
Tv8ny6XQLz9FibFqxSSq+1kOuJaDa7sNU7ExrzHqu6kYWTgVJGDBL4p88b00TYWb
aZ8f1ddklSGtItE+akzp885fNxemt64udgaMKYIMR1bbsqxfEz3ot3M+C2fezOCG
OHtlnm1aZ9miadRDNRT4V1jtW7YEzFrcV6Se6dPsckkHXE0XLQ4aujgJqJB9pRKx
luMTDPSigUPAebiB7bcKxKy3KhFuVNHmGDPqqdC+7mZ963Gmnmq9xx+89VhuK16z
tP857YI6Q3mJyPhB5TkzUjpRjhf+ML2wmER8PRvdvHrDXtaqaVrxyTt/Y0Sgn0N8
nQjfPmUsBMfloXZ86CESV+hZ4Da8/hTKRUicGjfAIUsmck/uBQMgSPXflKLTyoWe
u13MTXlk6IHlRrwBaZN81m56+yiEaob9truZgsxiu+FOQIs5LNmErySYjJeDEHAm
BLE7GOYhXNHYIvsj+vZGzJtGh3B4QoUT2BAVUGlzFn1vqz0McCj9DFGVXXeZ9P8A
OJ4ceMgOcwOhhcGDPJj6CgoismJx6J0wiVJsd0768WxPvBDzNN0sA0QVnUHZ5RpL
O8JJPo0UwREP3AMFnYswrFf9Rw5b6hUeIdr5OeiKMSXGHjBFXceTCDMLdQnrfzX/
Snnb8zMvK4wweSkmZi+WWdzavqk8OeENG1wU+mji1eUBTJ0aLqHhMqJiavenGaet
nc1HNskRhF33xOkCWF1UVHEJ94615GeUbrIzIYFRwTGkWAKxxnKk9xxeIx90NDzG
mN/dNNmOQEP7jmQxWWpUTIK7YHOw/7HlFzYnHzOHSZIGXCH6Yr+7wosR4WfOayXq
fkawNFKwqPATYfvKJd7j3QnNta0aKYnwvq4nGO8rjmfpzq66MTXNosAnEW/1/YXw
ghugANKto3oY0wIgDMCGDUYBo5fJ3lnaYhpTZOuDM5KcOHETf5i650stzKxAQuaq
95hTyj4q8en+Pypn5tI50dohbC4S1ogFmg3o3Dkm5I4pMGYLB7nHxeHbbC22cpsa
AUjaj/74zmqo6iq4j4AWVxcj9Jpsl1dU11r5oDO032QUwvPiDmUfVNM+FLRtynyc
VRPvHYU9n9iysQlEoy5E1eHa/sOuhrU0+mwWh8mfBNL8SIJViEBZClLmLAnPwM/N
BR8PEyBMqExIxcFcFvgh1rkqS4vug5A2ixVdC21eCbv2utTQlyxj2URWTiVfmZkm
Gy/uzo9jg+YbO2RBFsY7l7vO/acDJ3YR/xAmo23BHqQmpgdnVnWkymLZ5whvvSnW
NnKJ0YMPw5AuLY1nrf9d8MB0GhwoIPlC60hNyL7+Hr7AWvcGF+6fnkltmqWsoQEG
L0CCxhfjg6F69bgHdJ9tF9mB+gOiknU/rJkb1a2ym3W9V+wgtmJiGh/Il+sGEsH2
NksHGxMJiaGuW9zlDIZTw6zTxLCoVhB0grvPqvaeRPkLrwEQH0sGT1AciGtY/n8E
7BYhIdssqpvEWZW1AD3LWz9LK8khVmvbqNiBq1f6sImnjs1xyRQMSEVt8WCIxuCo
uYGsipwzUIWNKI4fiiIyIwPcC/DNfHktofVJWRDiSp9fuummEwKXT/NJDfzsTo7N
UaZs0IZIlyS/vUwcqrNy+qs/PXeEwqYSilyDa+GU8ZqPXIIp1lwFxzNqEGGOUBUN
fgj4PRG8pQzVLzmoEykHQLS0Xh/yoX2MrrGX/sDMRf2eMAN36FCIZeBCHW3HXvf2
KmJFAqFhRnzbeGQ/gE9++ekMYu4T0RUomfcfIrWI5198Mx6IB8dPULuw2A0MyfuY
3LosrKFkuFi4UDOluwvKmYx4iIeoh8Q/JyArSZzH0gUBxOHdpcys+L/hOsaIXOT/
v97QgH4TpoqTyY98TcOvBLFzRizLos0usVywTGKu0B9v4gyB3DpPDe+OmCGVHIN1
7rDenEf0rsItduezl2Aq/VCP87tI31mIUXVeX1nQSqW3/+J2OD5voTdgxzn5t3LV
N9UkQ+2xgX79spzfkDSv6fKkOQwpQPDgw9MJjCpJhDS+4pDYqi16ECpAtfcPywfU
8EShR3HCxDnyF2tAdYb9wQ==
`pragma protect end_protected
