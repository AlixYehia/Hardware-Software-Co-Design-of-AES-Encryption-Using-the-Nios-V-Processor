// AES_encrypt.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module AES_encrypt (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] intel_niosv_m_0_data_manager_awaddr;                            // intel_niosv_m_0:data_manager_awaddr -> mm_interconnect_0:intel_niosv_m_0_data_manager_awaddr
	wire   [1:0] intel_niosv_m_0_data_manager_bresp;                             // mm_interconnect_0:intel_niosv_m_0_data_manager_bresp -> intel_niosv_m_0:data_manager_bresp
	wire         intel_niosv_m_0_data_manager_arready;                           // mm_interconnect_0:intel_niosv_m_0_data_manager_arready -> intel_niosv_m_0:data_manager_arready
	wire  [31:0] intel_niosv_m_0_data_manager_rdata;                             // mm_interconnect_0:intel_niosv_m_0_data_manager_rdata -> intel_niosv_m_0:data_manager_rdata
	wire   [3:0] intel_niosv_m_0_data_manager_wstrb;                             // intel_niosv_m_0:data_manager_wstrb -> mm_interconnect_0:intel_niosv_m_0_data_manager_wstrb
	wire         intel_niosv_m_0_data_manager_wready;                            // mm_interconnect_0:intel_niosv_m_0_data_manager_wready -> intel_niosv_m_0:data_manager_wready
	wire         intel_niosv_m_0_data_manager_awready;                           // mm_interconnect_0:intel_niosv_m_0_data_manager_awready -> intel_niosv_m_0:data_manager_awready
	wire         intel_niosv_m_0_data_manager_rready;                            // intel_niosv_m_0:data_manager_rready -> mm_interconnect_0:intel_niosv_m_0_data_manager_rready
	wire         intel_niosv_m_0_data_manager_bready;                            // intel_niosv_m_0:data_manager_bready -> mm_interconnect_0:intel_niosv_m_0_data_manager_bready
	wire         intel_niosv_m_0_data_manager_wvalid;                            // intel_niosv_m_0:data_manager_wvalid -> mm_interconnect_0:intel_niosv_m_0_data_manager_wvalid
	wire  [31:0] intel_niosv_m_0_data_manager_araddr;                            // intel_niosv_m_0:data_manager_araddr -> mm_interconnect_0:intel_niosv_m_0_data_manager_araddr
	wire   [2:0] intel_niosv_m_0_data_manager_arprot;                            // intel_niosv_m_0:data_manager_arprot -> mm_interconnect_0:intel_niosv_m_0_data_manager_arprot
	wire   [1:0] intel_niosv_m_0_data_manager_rresp;                             // mm_interconnect_0:intel_niosv_m_0_data_manager_rresp -> intel_niosv_m_0:data_manager_rresp
	wire   [2:0] intel_niosv_m_0_data_manager_awprot;                            // intel_niosv_m_0:data_manager_awprot -> mm_interconnect_0:intel_niosv_m_0_data_manager_awprot
	wire  [31:0] intel_niosv_m_0_data_manager_wdata;                             // intel_niosv_m_0:data_manager_wdata -> mm_interconnect_0:intel_niosv_m_0_data_manager_wdata
	wire         intel_niosv_m_0_data_manager_arvalid;                           // intel_niosv_m_0:data_manager_arvalid -> mm_interconnect_0:intel_niosv_m_0_data_manager_arvalid
	wire         intel_niosv_m_0_data_manager_bvalid;                            // mm_interconnect_0:intel_niosv_m_0_data_manager_bvalid -> intel_niosv_m_0:data_manager_bvalid
	wire         intel_niosv_m_0_data_manager_awvalid;                           // intel_niosv_m_0:data_manager_awvalid -> mm_interconnect_0:intel_niosv_m_0_data_manager_awvalid
	wire         intel_niosv_m_0_data_manager_rvalid;                            // mm_interconnect_0:intel_niosv_m_0_data_manager_rvalid -> intel_niosv_m_0:data_manager_rvalid
	wire  [31:0] intel_niosv_m_0_instruction_manager_awaddr;                     // intel_niosv_m_0:instruction_manager_awaddr -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_awaddr
	wire   [1:0] intel_niosv_m_0_instruction_manager_bresp;                      // mm_interconnect_0:intel_niosv_m_0_instruction_manager_bresp -> intel_niosv_m_0:instruction_manager_bresp
	wire         intel_niosv_m_0_instruction_manager_arready;                    // mm_interconnect_0:intel_niosv_m_0_instruction_manager_arready -> intel_niosv_m_0:instruction_manager_arready
	wire  [31:0] intel_niosv_m_0_instruction_manager_rdata;                      // mm_interconnect_0:intel_niosv_m_0_instruction_manager_rdata -> intel_niosv_m_0:instruction_manager_rdata
	wire   [3:0] intel_niosv_m_0_instruction_manager_wstrb;                      // intel_niosv_m_0:instruction_manager_wstrb -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_wstrb
	wire         intel_niosv_m_0_instruction_manager_wready;                     // mm_interconnect_0:intel_niosv_m_0_instruction_manager_wready -> intel_niosv_m_0:instruction_manager_wready
	wire         intel_niosv_m_0_instruction_manager_awready;                    // mm_interconnect_0:intel_niosv_m_0_instruction_manager_awready -> intel_niosv_m_0:instruction_manager_awready
	wire         intel_niosv_m_0_instruction_manager_rready;                     // intel_niosv_m_0:instruction_manager_rready -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_rready
	wire         intel_niosv_m_0_instruction_manager_bready;                     // intel_niosv_m_0:instruction_manager_bready -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_bready
	wire         intel_niosv_m_0_instruction_manager_wvalid;                     // intel_niosv_m_0:instruction_manager_wvalid -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_wvalid
	wire  [31:0] intel_niosv_m_0_instruction_manager_araddr;                     // intel_niosv_m_0:instruction_manager_araddr -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_araddr
	wire   [2:0] intel_niosv_m_0_instruction_manager_arprot;                     // intel_niosv_m_0:instruction_manager_arprot -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_arprot
	wire   [1:0] intel_niosv_m_0_instruction_manager_rresp;                      // mm_interconnect_0:intel_niosv_m_0_instruction_manager_rresp -> intel_niosv_m_0:instruction_manager_rresp
	wire   [2:0] intel_niosv_m_0_instruction_manager_awprot;                     // intel_niosv_m_0:instruction_manager_awprot -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_awprot
	wire  [31:0] intel_niosv_m_0_instruction_manager_wdata;                      // intel_niosv_m_0:instruction_manager_wdata -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_wdata
	wire         intel_niosv_m_0_instruction_manager_arvalid;                    // intel_niosv_m_0:instruction_manager_arvalid -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_arvalid
	wire         intel_niosv_m_0_instruction_manager_bvalid;                     // mm_interconnect_0:intel_niosv_m_0_instruction_manager_bvalid -> intel_niosv_m_0:instruction_manager_bvalid
	wire         intel_niosv_m_0_instruction_manager_awvalid;                    // intel_niosv_m_0:instruction_manager_awvalid -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_awvalid
	wire         intel_niosv_m_0_instruction_manager_rvalid;                     // mm_interconnect_0:intel_niosv_m_0_instruction_manager_rvalid -> intel_niosv_m_0:instruction_manager_rvalid
	wire   [5:0] mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_awaddr;       // mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_awaddr -> AES_AXI_0:S_AXI_AWADDR
	wire   [1:0] mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_bresp;        // AES_AXI_0:S_AXI_BRESP -> mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_bresp
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_arready;      // AES_AXI_0:S_AXI_ARREADY -> mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_arready
	wire  [31:0] mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rdata;        // AES_AXI_0:S_AXI_RDATA -> mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_rdata
	wire   [3:0] mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wstrb;        // mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_wstrb -> AES_AXI_0:S_AXI_WSTRB
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wready;       // AES_AXI_0:S_AXI_WREADY -> mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_wready
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_awready;      // AES_AXI_0:S_AXI_AWREADY -> mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_awready
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rready;       // mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_rready -> AES_AXI_0:S_AXI_RREADY
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_bready;       // mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_bready -> AES_AXI_0:S_AXI_BREADY
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wvalid;       // mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_wvalid -> AES_AXI_0:S_AXI_WVALID
	wire   [5:0] mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_araddr;       // mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_araddr -> AES_AXI_0:S_AXI_ARADDR
	wire   [1:0] mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rresp;        // AES_AXI_0:S_AXI_RRESP -> mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_rresp
	wire  [31:0] mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wdata;        // mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_wdata -> AES_AXI_0:S_AXI_WDATA
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_arvalid;      // mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_arvalid -> AES_AXI_0:S_AXI_ARVALID
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_bvalid;       // AES_AXI_0:S_AXI_BVALID -> mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_bvalid
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_awvalid;      // mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_awvalid -> AES_AXI_0:S_AXI_AWVALID
	wire         mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rvalid;       // AES_AXI_0:S_AXI_RVALID -> mm_interconnect_0:AES_AXI_0_altera_axi4lite_slave_rvalid
	wire   [5:0] mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_awaddr;      // mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_awaddr -> AES_DECR_0:S_AXI_AWADDR
	wire   [1:0] mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_bresp;       // AES_DECR_0:S_AXI_BRESP -> mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_bresp
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_arready;     // AES_DECR_0:S_AXI_ARREADY -> mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_arready
	wire  [31:0] mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rdata;       // AES_DECR_0:S_AXI_RDATA -> mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_rdata
	wire   [3:0] mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wstrb;       // mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_wstrb -> AES_DECR_0:S_AXI_WSTRB
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wready;      // AES_DECR_0:S_AXI_WREADY -> mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_wready
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_awready;     // AES_DECR_0:S_AXI_AWREADY -> mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_awready
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rready;      // mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_rready -> AES_DECR_0:S_AXI_RREADY
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_bready;      // mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_bready -> AES_DECR_0:S_AXI_BREADY
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wvalid;      // mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_wvalid -> AES_DECR_0:S_AXI_WVALID
	wire   [5:0] mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_araddr;      // mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_araddr -> AES_DECR_0:S_AXI_ARADDR
	wire   [1:0] mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rresp;       // AES_DECR_0:S_AXI_RRESP -> mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_rresp
	wire  [31:0] mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wdata;       // mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_wdata -> AES_DECR_0:S_AXI_WDATA
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_arvalid;     // mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_arvalid -> AES_DECR_0:S_AXI_ARVALID
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_bvalid;      // AES_DECR_0:S_AXI_BVALID -> mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_bvalid
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_awvalid;     // mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_awvalid -> AES_DECR_0:S_AXI_AWVALID
	wire         mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rvalid;      // AES_DECR_0:S_AXI_RVALID -> mm_interconnect_0:AES_DECR_0_altera_axi4lite_slave_rvalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;       // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;    // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata;            // intel_niosv_m_0:dm_agent_readdata -> mm_interconnect_0:intel_niosv_m_0_dm_agent_readdata
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest;         // intel_niosv_m_0:dm_agent_waitrequest -> mm_interconnect_0:intel_niosv_m_0_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_address;             // mm_interconnect_0:intel_niosv_m_0_dm_agent_address -> intel_niosv_m_0:dm_agent_address
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_read;                // mm_interconnect_0:intel_niosv_m_0_dm_agent_read -> intel_niosv_m_0:dm_agent_read
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid;       // intel_niosv_m_0:dm_agent_readdatavalid -> mm_interconnect_0:intel_niosv_m_0_dm_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_write;               // mm_interconnect_0:intel_niosv_m_0_dm_agent_write -> intel_niosv_m_0:dm_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata;           // mm_interconnect_0:intel_niosv_m_0_dm_agent_writedata -> intel_niosv_m_0:dm_agent_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;               // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                 // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_0_s1_address;                  // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;               // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                    // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                    // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata;      // intel_niosv_m_0:timer_sw_agent_readdata -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_readdata
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest;   // intel_niosv_m_0:timer_sw_agent_waitrequest -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address;       // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_address -> intel_niosv_m_0:timer_sw_agent_address
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read;          // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_read -> intel_niosv_m_0:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable;    // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_byteenable -> intel_niosv_m_0:timer_sw_agent_byteenable
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid; // intel_niosv_m_0:timer_sw_agent_readdatavalid -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write;         // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_write -> intel_niosv_m_0:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata;     // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_writedata -> intel_niosv_m_0:timer_sw_agent_writedata
	wire         irq_mapper_receiver0_irq;                                       // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [15:0] intel_niosv_m_0_platform_irq_rx_irq;                            // irq_mapper:sender_irq -> intel_niosv_m_0:platform_irq_rx_irq
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [AES_AXI_0:ARESETN, AES_DECR_0:ARESETN, intel_niosv_m_0:reset_reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:intel_niosv_m_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                             // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	AES_AXI_wrapper #(
		.ADDR_WIDTH (6),
		.DATA_WIDTH (32)
	) aes_axi_0 (
		.ACLK          (clk_clk),                                                   //            clock_sink.clk
		.ARESETN       (~rst_controller_reset_out_reset),                           //            reset_sink.reset_n
		.S_AXI_AWADDR  (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_awaddr),  // altera_axi4lite_slave.awaddr
		.S_AXI_AWVALID (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_awvalid), //                      .awvalid
		.S_AXI_AWREADY (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_awready), //                      .awready
		.S_AXI_WDATA   (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wdata),   //                      .wdata
		.S_AXI_WSTRB   (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wstrb),   //                      .wstrb
		.S_AXI_WVALID  (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wvalid),  //                      .wvalid
		.S_AXI_WREADY  (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wready),  //                      .wready
		.S_AXI_BRESP   (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_bresp),   //                      .bresp
		.S_AXI_BVALID  (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_bvalid),  //                      .bvalid
		.S_AXI_BREADY  (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_bready),  //                      .bready
		.S_AXI_ARADDR  (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_araddr),  //                      .araddr
		.S_AXI_ARVALID (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_arvalid), //                      .arvalid
		.S_AXI_ARREADY (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_arready), //                      .arready
		.S_AXI_RDATA   (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rdata),   //                      .rdata
		.S_AXI_RRESP   (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rresp),   //                      .rresp
		.S_AXI_RVALID  (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rvalid),  //                      .rvalid
		.S_AXI_RREADY  (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rready)   //                      .rready
	);

	AES_DEC_AXI_wrapper #(
		.ADDR_WIDTH (6),
		.DATA_WIDTH (32)
	) aes_decr_0 (
		.ACLK          (clk_clk),                                                    //            clock_sink.clk
		.ARESETN       (~rst_controller_reset_out_reset),                            //            reset_sink.reset_n
		.S_AXI_AWADDR  (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_awaddr),  // altera_axi4lite_slave.awaddr
		.S_AXI_AWVALID (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_awvalid), //                      .awvalid
		.S_AXI_AWREADY (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_awready), //                      .awready
		.S_AXI_WDATA   (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wdata),   //                      .wdata
		.S_AXI_WSTRB   (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wstrb),   //                      .wstrb
		.S_AXI_WVALID  (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wvalid),  //                      .wvalid
		.S_AXI_WREADY  (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wready),  //                      .wready
		.S_AXI_BRESP   (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_bresp),   //                      .bresp
		.S_AXI_BVALID  (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_bvalid),  //                      .bvalid
		.S_AXI_BREADY  (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_bready),  //                      .bready
		.S_AXI_ARADDR  (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_araddr),  //                      .araddr
		.S_AXI_ARVALID (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_arvalid), //                      .arvalid
		.S_AXI_ARREADY (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_arready), //                      .arready
		.S_AXI_RDATA   (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rdata),   //                      .rdata
		.S_AXI_RRESP   (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rresp),   //                      .rresp
		.S_AXI_RVALID  (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rvalid),  //                      .rvalid
		.S_AXI_RREADY  (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rready)   //                      .rready
	);

	AES_encrypt_intel_niosv_m_0 intel_niosv_m_0 (
		.clk                          (clk_clk),                                                        //                 clk.clk
		.reset_reset                  (rst_controller_reset_out_reset),                                 //               reset.reset
		.platform_irq_rx_irq          (intel_niosv_m_0_platform_irq_rx_irq),                            //     platform_irq_rx.irq
		.timer_sw_agent_address       (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address),       //      timer_sw_agent.address
		.timer_sw_agent_byteenable    (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable),    //                    .byteenable
		.timer_sw_agent_read          (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read),          //                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata),      //                    .readdata
		.timer_sw_agent_write         (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write),         //                    .write
		.timer_sw_agent_writedata     (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata),     //                    .writedata
		.timer_sw_agent_waitrequest   (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest),   //                    .waitrequest
		.timer_sw_agent_readdatavalid (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid), //                    .readdatavalid
		.instruction_manager_awaddr   (intel_niosv_m_0_instruction_manager_awaddr),                     // instruction_manager.awaddr
		.instruction_manager_awprot   (intel_niosv_m_0_instruction_manager_awprot),                     //                    .awprot
		.instruction_manager_awvalid  (intel_niosv_m_0_instruction_manager_awvalid),                    //                    .awvalid
		.instruction_manager_awready  (intel_niosv_m_0_instruction_manager_awready),                    //                    .awready
		.instruction_manager_wdata    (intel_niosv_m_0_instruction_manager_wdata),                      //                    .wdata
		.instruction_manager_wstrb    (intel_niosv_m_0_instruction_manager_wstrb),                      //                    .wstrb
		.instruction_manager_wvalid   (intel_niosv_m_0_instruction_manager_wvalid),                     //                    .wvalid
		.instruction_manager_wready   (intel_niosv_m_0_instruction_manager_wready),                     //                    .wready
		.instruction_manager_bresp    (intel_niosv_m_0_instruction_manager_bresp),                      //                    .bresp
		.instruction_manager_bvalid   (intel_niosv_m_0_instruction_manager_bvalid),                     //                    .bvalid
		.instruction_manager_bready   (intel_niosv_m_0_instruction_manager_bready),                     //                    .bready
		.instruction_manager_araddr   (intel_niosv_m_0_instruction_manager_araddr),                     //                    .araddr
		.instruction_manager_arprot   (intel_niosv_m_0_instruction_manager_arprot),                     //                    .arprot
		.instruction_manager_arvalid  (intel_niosv_m_0_instruction_manager_arvalid),                    //                    .arvalid
		.instruction_manager_arready  (intel_niosv_m_0_instruction_manager_arready),                    //                    .arready
		.instruction_manager_rdata    (intel_niosv_m_0_instruction_manager_rdata),                      //                    .rdata
		.instruction_manager_rresp    (intel_niosv_m_0_instruction_manager_rresp),                      //                    .rresp
		.instruction_manager_rvalid   (intel_niosv_m_0_instruction_manager_rvalid),                     //                    .rvalid
		.instruction_manager_rready   (intel_niosv_m_0_instruction_manager_rready),                     //                    .rready
		.data_manager_awaddr          (intel_niosv_m_0_data_manager_awaddr),                            //        data_manager.awaddr
		.data_manager_awprot          (intel_niosv_m_0_data_manager_awprot),                            //                    .awprot
		.data_manager_awvalid         (intel_niosv_m_0_data_manager_awvalid),                           //                    .awvalid
		.data_manager_awready         (intel_niosv_m_0_data_manager_awready),                           //                    .awready
		.data_manager_wdata           (intel_niosv_m_0_data_manager_wdata),                             //                    .wdata
		.data_manager_wstrb           (intel_niosv_m_0_data_manager_wstrb),                             //                    .wstrb
		.data_manager_wvalid          (intel_niosv_m_0_data_manager_wvalid),                            //                    .wvalid
		.data_manager_wready          (intel_niosv_m_0_data_manager_wready),                            //                    .wready
		.data_manager_bresp           (intel_niosv_m_0_data_manager_bresp),                             //                    .bresp
		.data_manager_bvalid          (intel_niosv_m_0_data_manager_bvalid),                            //                    .bvalid
		.data_manager_bready          (intel_niosv_m_0_data_manager_bready),                            //                    .bready
		.data_manager_araddr          (intel_niosv_m_0_data_manager_araddr),                            //                    .araddr
		.data_manager_arprot          (intel_niosv_m_0_data_manager_arprot),                            //                    .arprot
		.data_manager_arvalid         (intel_niosv_m_0_data_manager_arvalid),                           //                    .arvalid
		.data_manager_arready         (intel_niosv_m_0_data_manager_arready),                           //                    .arready
		.data_manager_rdata           (intel_niosv_m_0_data_manager_rdata),                             //                    .rdata
		.data_manager_rresp           (intel_niosv_m_0_data_manager_rresp),                             //                    .rresp
		.data_manager_rvalid          (intel_niosv_m_0_data_manager_rvalid),                            //                    .rvalid
		.data_manager_rready          (intel_niosv_m_0_data_manager_rready),                            //                    .rready
		.dm_agent_address             (mm_interconnect_0_intel_niosv_m_0_dm_agent_address),             //            dm_agent.address
		.dm_agent_read                (mm_interconnect_0_intel_niosv_m_0_dm_agent_read),                //                    .read
		.dm_agent_readdata            (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata),            //                    .readdata
		.dm_agent_write               (mm_interconnect_0_intel_niosv_m_0_dm_agent_write),               //                    .write
		.dm_agent_writedata           (mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata),           //                    .writedata
		.dm_agent_waitrequest         (mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest),         //                    .waitrequest
		.dm_agent_readdatavalid       (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid)        //                    .readdatavalid
	);

	altera_avalon_jtag_uart #(
		.readBufferDepth            (32),
		.readIRQThreshold           (8),
		.useRegistersForReadBuffer  (0),
		.useRegistersForWriteBuffer (0),
		.writeBufferDepth           (32),
		.writeIRQThreshold          (8),
		.printingMethod             (0),
		.FIFO_WIDTH                 (8),
		.WR_WIDTHU                  (5),
		.RD_WIDTHU                  (5),
		.write_le                   ("ON"),
		.read_le                    ("ON"),
		.HEX_WRITE_DEPTH_STR        (32),
		.HEX_READ_DEPTH_STR         (32),
		.legacySignalAllow          (0)
	) jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	AES_encrypt_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	AES_encrypt_mm_interconnect_0 mm_interconnect_0 (
		.AES_AXI_0_altera_axi4lite_slave_awaddr            (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_awaddr),       //             AES_AXI_0_altera_axi4lite_slave.awaddr
		.AES_AXI_0_altera_axi4lite_slave_awprot            (),                                                               //                                            .awprot
		.AES_AXI_0_altera_axi4lite_slave_awvalid           (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_awvalid),      //                                            .awvalid
		.AES_AXI_0_altera_axi4lite_slave_awready           (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_awready),      //                                            .awready
		.AES_AXI_0_altera_axi4lite_slave_wdata             (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wdata),        //                                            .wdata
		.AES_AXI_0_altera_axi4lite_slave_wstrb             (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wstrb),        //                                            .wstrb
		.AES_AXI_0_altera_axi4lite_slave_wvalid            (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wvalid),       //                                            .wvalid
		.AES_AXI_0_altera_axi4lite_slave_wready            (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_wready),       //                                            .wready
		.AES_AXI_0_altera_axi4lite_slave_bresp             (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_bresp),        //                                            .bresp
		.AES_AXI_0_altera_axi4lite_slave_bvalid            (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_bvalid),       //                                            .bvalid
		.AES_AXI_0_altera_axi4lite_slave_bready            (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_bready),       //                                            .bready
		.AES_AXI_0_altera_axi4lite_slave_araddr            (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_araddr),       //                                            .araddr
		.AES_AXI_0_altera_axi4lite_slave_arprot            (),                                                               //                                            .arprot
		.AES_AXI_0_altera_axi4lite_slave_arvalid           (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_arvalid),      //                                            .arvalid
		.AES_AXI_0_altera_axi4lite_slave_arready           (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_arready),      //                                            .arready
		.AES_AXI_0_altera_axi4lite_slave_rdata             (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rdata),        //                                            .rdata
		.AES_AXI_0_altera_axi4lite_slave_rresp             (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rresp),        //                                            .rresp
		.AES_AXI_0_altera_axi4lite_slave_rvalid            (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rvalid),       //                                            .rvalid
		.AES_AXI_0_altera_axi4lite_slave_rready            (mm_interconnect_0_aes_axi_0_altera_axi4lite_slave_rready),       //                                            .rready
		.AES_DECR_0_altera_axi4lite_slave_awaddr           (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_awaddr),      //            AES_DECR_0_altera_axi4lite_slave.awaddr
		.AES_DECR_0_altera_axi4lite_slave_awprot           (),                                                               //                                            .awprot
		.AES_DECR_0_altera_axi4lite_slave_awvalid          (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_awvalid),     //                                            .awvalid
		.AES_DECR_0_altera_axi4lite_slave_awready          (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_awready),     //                                            .awready
		.AES_DECR_0_altera_axi4lite_slave_wdata            (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wdata),       //                                            .wdata
		.AES_DECR_0_altera_axi4lite_slave_wstrb            (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wstrb),       //                                            .wstrb
		.AES_DECR_0_altera_axi4lite_slave_wvalid           (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wvalid),      //                                            .wvalid
		.AES_DECR_0_altera_axi4lite_slave_wready           (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_wready),      //                                            .wready
		.AES_DECR_0_altera_axi4lite_slave_bresp            (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_bresp),       //                                            .bresp
		.AES_DECR_0_altera_axi4lite_slave_bvalid           (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_bvalid),      //                                            .bvalid
		.AES_DECR_0_altera_axi4lite_slave_bready           (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_bready),      //                                            .bready
		.AES_DECR_0_altera_axi4lite_slave_araddr           (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_araddr),      //                                            .araddr
		.AES_DECR_0_altera_axi4lite_slave_arprot           (),                                                               //                                            .arprot
		.AES_DECR_0_altera_axi4lite_slave_arvalid          (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_arvalid),     //                                            .arvalid
		.AES_DECR_0_altera_axi4lite_slave_arready          (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_arready),     //                                            .arready
		.AES_DECR_0_altera_axi4lite_slave_rdata            (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rdata),       //                                            .rdata
		.AES_DECR_0_altera_axi4lite_slave_rresp            (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rresp),       //                                            .rresp
		.AES_DECR_0_altera_axi4lite_slave_rvalid           (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rvalid),      //                                            .rvalid
		.AES_DECR_0_altera_axi4lite_slave_rready           (mm_interconnect_0_aes_decr_0_altera_axi4lite_slave_rready),      //                                            .rready
		.intel_niosv_m_0_data_manager_awaddr               (intel_niosv_m_0_data_manager_awaddr),                            //                intel_niosv_m_0_data_manager.awaddr
		.intel_niosv_m_0_data_manager_awprot               (intel_niosv_m_0_data_manager_awprot),                            //                                            .awprot
		.intel_niosv_m_0_data_manager_awvalid              (intel_niosv_m_0_data_manager_awvalid),                           //                                            .awvalid
		.intel_niosv_m_0_data_manager_awready              (intel_niosv_m_0_data_manager_awready),                           //                                            .awready
		.intel_niosv_m_0_data_manager_wdata                (intel_niosv_m_0_data_manager_wdata),                             //                                            .wdata
		.intel_niosv_m_0_data_manager_wstrb                (intel_niosv_m_0_data_manager_wstrb),                             //                                            .wstrb
		.intel_niosv_m_0_data_manager_wvalid               (intel_niosv_m_0_data_manager_wvalid),                            //                                            .wvalid
		.intel_niosv_m_0_data_manager_wready               (intel_niosv_m_0_data_manager_wready),                            //                                            .wready
		.intel_niosv_m_0_data_manager_bresp                (intel_niosv_m_0_data_manager_bresp),                             //                                            .bresp
		.intel_niosv_m_0_data_manager_bvalid               (intel_niosv_m_0_data_manager_bvalid),                            //                                            .bvalid
		.intel_niosv_m_0_data_manager_bready               (intel_niosv_m_0_data_manager_bready),                            //                                            .bready
		.intel_niosv_m_0_data_manager_araddr               (intel_niosv_m_0_data_manager_araddr),                            //                                            .araddr
		.intel_niosv_m_0_data_manager_arprot               (intel_niosv_m_0_data_manager_arprot),                            //                                            .arprot
		.intel_niosv_m_0_data_manager_arvalid              (intel_niosv_m_0_data_manager_arvalid),                           //                                            .arvalid
		.intel_niosv_m_0_data_manager_arready              (intel_niosv_m_0_data_manager_arready),                           //                                            .arready
		.intel_niosv_m_0_data_manager_rdata                (intel_niosv_m_0_data_manager_rdata),                             //                                            .rdata
		.intel_niosv_m_0_data_manager_rresp                (intel_niosv_m_0_data_manager_rresp),                             //                                            .rresp
		.intel_niosv_m_0_data_manager_rvalid               (intel_niosv_m_0_data_manager_rvalid),                            //                                            .rvalid
		.intel_niosv_m_0_data_manager_rready               (intel_niosv_m_0_data_manager_rready),                            //                                            .rready
		.intel_niosv_m_0_instruction_manager_awaddr        (intel_niosv_m_0_instruction_manager_awaddr),                     //         intel_niosv_m_0_instruction_manager.awaddr
		.intel_niosv_m_0_instruction_manager_awprot        (intel_niosv_m_0_instruction_manager_awprot),                     //                                            .awprot
		.intel_niosv_m_0_instruction_manager_awvalid       (intel_niosv_m_0_instruction_manager_awvalid),                    //                                            .awvalid
		.intel_niosv_m_0_instruction_manager_awready       (intel_niosv_m_0_instruction_manager_awready),                    //                                            .awready
		.intel_niosv_m_0_instruction_manager_wdata         (intel_niosv_m_0_instruction_manager_wdata),                      //                                            .wdata
		.intel_niosv_m_0_instruction_manager_wstrb         (intel_niosv_m_0_instruction_manager_wstrb),                      //                                            .wstrb
		.intel_niosv_m_0_instruction_manager_wvalid        (intel_niosv_m_0_instruction_manager_wvalid),                     //                                            .wvalid
		.intel_niosv_m_0_instruction_manager_wready        (intel_niosv_m_0_instruction_manager_wready),                     //                                            .wready
		.intel_niosv_m_0_instruction_manager_bresp         (intel_niosv_m_0_instruction_manager_bresp),                      //                                            .bresp
		.intel_niosv_m_0_instruction_manager_bvalid        (intel_niosv_m_0_instruction_manager_bvalid),                     //                                            .bvalid
		.intel_niosv_m_0_instruction_manager_bready        (intel_niosv_m_0_instruction_manager_bready),                     //                                            .bready
		.intel_niosv_m_0_instruction_manager_araddr        (intel_niosv_m_0_instruction_manager_araddr),                     //                                            .araddr
		.intel_niosv_m_0_instruction_manager_arprot        (intel_niosv_m_0_instruction_manager_arprot),                     //                                            .arprot
		.intel_niosv_m_0_instruction_manager_arvalid       (intel_niosv_m_0_instruction_manager_arvalid),                    //                                            .arvalid
		.intel_niosv_m_0_instruction_manager_arready       (intel_niosv_m_0_instruction_manager_arready),                    //                                            .arready
		.intel_niosv_m_0_instruction_manager_rdata         (intel_niosv_m_0_instruction_manager_rdata),                      //                                            .rdata
		.intel_niosv_m_0_instruction_manager_rresp         (intel_niosv_m_0_instruction_manager_rresp),                      //                                            .rresp
		.intel_niosv_m_0_instruction_manager_rvalid        (intel_niosv_m_0_instruction_manager_rvalid),                     //                                            .rvalid
		.intel_niosv_m_0_instruction_manager_rready        (intel_niosv_m_0_instruction_manager_rready),                     //                                            .rready
		.clk_0_clk_clk                                     (clk_clk),                                                        //                                   clk_0_clk.clk
		.intel_niosv_m_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // intel_niosv_m_0_reset_reset_bridge_in_reset.reset
		.intel_niosv_m_0_dm_agent_address                  (mm_interconnect_0_intel_niosv_m_0_dm_agent_address),             //                    intel_niosv_m_0_dm_agent.address
		.intel_niosv_m_0_dm_agent_write                    (mm_interconnect_0_intel_niosv_m_0_dm_agent_write),               //                                            .write
		.intel_niosv_m_0_dm_agent_read                     (mm_interconnect_0_intel_niosv_m_0_dm_agent_read),                //                                            .read
		.intel_niosv_m_0_dm_agent_readdata                 (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata),            //                                            .readdata
		.intel_niosv_m_0_dm_agent_writedata                (mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata),           //                                            .writedata
		.intel_niosv_m_0_dm_agent_readdatavalid            (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid),       //                                            .readdatavalid
		.intel_niosv_m_0_dm_agent_waitrequest              (mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest),         //                                            .waitrequest
		.intel_niosv_m_0_timer_sw_agent_address            (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address),       //              intel_niosv_m_0_timer_sw_agent.address
		.intel_niosv_m_0_timer_sw_agent_write              (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write),         //                                            .write
		.intel_niosv_m_0_timer_sw_agent_read               (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read),          //                                            .read
		.intel_niosv_m_0_timer_sw_agent_readdata           (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata),      //                                            .readdata
		.intel_niosv_m_0_timer_sw_agent_writedata          (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata),     //                                            .writedata
		.intel_niosv_m_0_timer_sw_agent_byteenable         (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable),    //                                            .byteenable
		.intel_niosv_m_0_timer_sw_agent_readdatavalid      (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid), //                                            .readdatavalid
		.intel_niosv_m_0_timer_sw_agent_waitrequest        (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest),   //                                            .waitrequest
		.jtag_uart_0_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),        //               jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),          //                                            .write
		.jtag_uart_0_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),           //                                            .read
		.jtag_uart_0_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),       //                                            .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),      //                                            .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),    //                                            .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),     //                                            .chipselect
		.onchip_memory2_0_s1_address                       (mm_interconnect_0_onchip_memory2_0_s1_address),                  //                         onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                         (mm_interconnect_0_onchip_memory2_0_s1_write),                    //                                            .write
		.onchip_memory2_0_s1_readdata                      (mm_interconnect_0_onchip_memory2_0_s1_readdata),                 //                                            .readdata
		.onchip_memory2_0_s1_writedata                     (mm_interconnect_0_onchip_memory2_0_s1_writedata),                //                                            .writedata
		.onchip_memory2_0_s1_byteenable                    (mm_interconnect_0_onchip_memory2_0_s1_byteenable),               //                                            .byteenable
		.onchip_memory2_0_s1_chipselect                    (mm_interconnect_0_onchip_memory2_0_s1_chipselect),               //                                            .chipselect
		.onchip_memory2_0_s1_clken                         (mm_interconnect_0_onchip_memory2_0_s1_clken)                     //                                            .clken
	);

	AES_encrypt_irq_mapper irq_mapper (
		.clk           (clk_clk),                             //       clk.clk
		.reset         (rst_controller_reset_out_reset),      // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),            // receiver0.irq
		.sender_irq    (intel_niosv_m_0_platform_irq_rx_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
