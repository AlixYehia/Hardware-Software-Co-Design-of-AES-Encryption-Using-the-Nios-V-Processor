// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
TbpdsbkTv9BOA7IBGsIpYM9sAhERJqMDuH9NNZ/M6moBXMcGoBX9qwM2br1JnoVp2guAyPIcdCrk
q35fPWaLcBPkLIH907zdaeMDyNYEkgIGawcWw7IOMKVnIZFso9D7heaxIRJllE5T0qj5uOJQd4i4
N+0EKZ/RcknKdnXPqanQiMosXVnyyDwsSznez3XfyZ8xudUFOfjDUrbxZMdkYAfc/vqrZ5jDHeKU
32r3UafYUvScuZOaLr3HPPqTjxK0qB53Z6M/q9vn9Mwv3I5OMg8nFzYXEL7S9AXEdPcCvFN2pUg+
chPD9yMDJjusq4UWNg+U3g3a9sbs5CQ7v8IqBg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 69152)
wGh5E51b/8NFAQFx7xiZm4urcqC0gnJeOPaxtSrjF9JYzDBwPGaNykCxcq57UrTT9Tr6GascPQiI
JbFQznTw+LmQ1HqMNbW5A7LDwfy0Y/CQYpTT5Uh5JZ3G3CS4CjoaIgvzKU/3jOyy50x0ls2G92uY
gvLyUEFjODPbzmzBOM5+eu4vQeUSsoJvEL2xGYy4qjsJs+ZPrg1ZzBHbvH4W5rX9Nw3jXxazDCmD
dnEyhslp6G7DlkKsZrU7KjTYMb7UZzU3HqpmiHG4gH6aFOn9T+R/zF7jG0VqFomSpEKr/waz48Uq
9y2y5DoblUIzuFgbQEjbF8T7TKCLqEzwqXBhSlfqNhBKLkMvptbznHDlGAquaVSGqymEzUaU4Z6l
5jLbJw0aWJFS7hG/6zNbBvak+iUoCbUEoHjCxrzzEGG4gI2hvUGxob9JI61p1Ock6mR652BcLhe5
rEycdwDeeJrRw8VPeUal0p/pFgEZCmmXKJHF6bp7rkf7lrcSJ4xqoM57AnI6EwQOJZmRmCuG8s33
t0rFg/WPR+vh3LiatLcdHFKtFWWWifuR6ObvOzjXPONOn21lLAwPkGlRm24hXW8wk1tuHYFCQnQe
m686ZY6bHQDmmqFPghGr9tD8y+DjdHyy3PNylDAD4Xuq6HSlWpGNJuErfkeRzN+GpRo76XZHwCSl
O2P637rABrz6RMqGh2gpFT/1niYhz+tC3B+bdT1CO1PFDr5MXCVnnB9BZT1qc/NkIuEBEfVAfko0
Pj/36MS1nq99BznIO352FH6t6T9+a76ObzK0ZnHCfJZevwc9x60Rj6tAQMYhtBUGY92c4c9urVb7
CYKluwuARRn+5l0WEDvRPhURvqLyCbdjRZzx7KISfI98WbuGbN0cmLI2TmBd2Zyc1VQYBPahZeMB
otpBhm9uIg5jyiBowXQ6aQ4H/2z0jhgfN/n+ihpQDfBB0oaOPx8SZO6bSFd7Prg2P/qeFGXyd1Gg
5+AhCa6eidKpjMtEAI1vXEfxOyw2dtDX5ok4KreX3x+MVLIIYobjeOZyIlTep5aj/L00Ujf1eDFA
Zh/QJvtvE4GIuASpbU/yYtObQdmh789kiLuEhcu51sDoL40ntyW1I2sjJxLXhnw+Scgr6/H+qC1A
rK20F/HjtxfEwvdDY95E7De/zVDFF5XeKBu3haFlFELUw067EQbXWe1KrZsGvSW07ngX7Bd2mlgC
u0bS2IeckxwYOY/LriLbkuF2ZPhAI3G7qM56DGqqFgOmb7Vg+thuEyT8ujgiLS/i41oiw9Wxc3Nc
K1ZBhLeM5nhRhoJCTlJY9ofGh+pa/1YhTiLya9AxyNl+PKLF/93cGGySgvd56kPrTsSkCTapCMFU
uXmQ1dlvbcQLv3/WlcWOj6XGLt5cNG/jzSJZMdkFi6YljUIq9NlrRNxFKFLvKWtREab5U17HNihw
ZCfSkHtJFy6i9yq3czmYRQTkEkNLMY0S1odIwnzCboV9yYyCmjaW6IAtz8ZRzcw1e/nwpYyJPVBA
rtYO8Hf7P5TX8syEvDoJecicTKNMhFL9jkiGCU58aaGa0aEqqjpAVtxnUav7bDRMABYZcBUyQ/pr
GlC1rH5317b0QiTnCzlqyWXtii5CDeUHff9iGkd+nzRv7GtGdlhtaU5bAF1UxMshDnhSrT7rH+F1
GW46sydMOtQekws8jMdW65V/QXQ94J0NJMbLnCVvhcCF5ADLtGRUUxWQcHkehxmAwWldys/Vn4Cr
1lujOCDHj6XMLgKpOkzkeQHMApmZzOCHzB2n+DM1rjfuKnKonqjS4dmiFF/SBjQABJUWPSriPYHi
j2pHozNoo2XXhC1TAOWPXjik9mI3NqrEqeMfodWlDuTQrg0EktET0VXkoZRgwspYbFqf0d1f4oJi
o4H6SkI5qPnMPW6vMBUf9UjtjGJTSjT6S9IdsNZcKxQw7Hay9QipUzipRsQhVO8oAEbwDIpRmfBb
feRgvcj9IiO+6UiYO7ZoQLOsf6NVOQPv22d4FiCBmlOBU6bqLE8sfCquRLHoHqU1nxnyDBPv11lB
/dsMpRZxV/BHmC8EGT3ZMdT85RIp6HGNvf8zQ7N9ZvXy2tb7HdcOlhWjvEfh0R/Ca1tJEtcMImqr
OE3PS5ItUnh2gecYFSGHlKC11NIvGSStA7NBJuUK16zTd2dRv5LZ1SuOoA4yxD6iy37R1ffuDeDQ
fiMMkDhEJm8lJzCeYBlDJDWQJ9GYWGkzvbBZrE3v8Vv+TKCG00m3WqSEanGcOPqzuJM/1feu02CD
l1Pps7rY2blm2/ldfY/bd+P5y6I6TTR00b32e/DCm2jnoELHWC0DvZK0wjYOraQCRqt1Dnf1nLLK
CU2fPqFhrIbQTLCcTK8yohikUllzQFjacHIsPuRjHfguxRxXUjSaY4R7tjUJAc3JlZcgVwMkP60+
LN7zbK4drPJ3uv7fLoGNBp0AmpDtSIAxwRmeD3dpKyTRwG5ycoWyLFoqmzdU3u36YFACgdkmgcBH
zbCqtn3U2I/HR7YiFV+SyEx+dTX8A8pp796BKDyjoJGjW7x0Gq0xH5DdK0+fEk0JSa5til6zcjIC
dDHjmTeZcej0OGnBP/eZfJzB7MZR1BfSBUfFSS/tdwcd3WbhS3aFH/0rsTlPcNrfyYE+HNEtMZhz
0ThJ44B5jgzrmViysL8+n1vVJc1Z487FxMYFJo+wpPwWGvVQBmxpsReYLIIh2Vab2sXb2l+DLrr6
HKTHA3e4K3MmT1eH0/VA/ZNckjSHz/CeVClKGFKPEHY21GsoZjR5+djqTVvRuAjuDenARLNfH9I8
3WTUewOsBV51IcryG04S86yBi48ePlML7qWUcEp75iSEdK85/aCmJ3EDwq++FRlXvj0jrQ3ZbwfR
ppSVAND57tgmd+D6Oal6sFkem446XTDv8lrvYek/y4wx3Uj3BcVA/kFhpZj+lf0O80+pYoUUVtA8
Q0HRvJZsJ5icTS3AM93yGw4USuLmkuODroRRJtf1T1cbdIgL5UNWbUyshEuSejj1Gx0dHcDlBeJO
FIuGoGoRZlNYXNoMht9v+BGIYAgJrBjRVT7bpYSPaKhOnWdpy5+N6UdKBIosEuLLrf+jpcVguNJf
ZUtUClE4/aWw75JFtakZySiWc9GFM43My+sTY5+odveemYRAnsh6z++6MmoAu0SC5n1qznhZ3qBD
l7XHow/6dupPeo/3yQwJxgwJMCc0i+IHrPChaq2f3pvmzcfKA0oSfwqvgWucc+t+tqC80+PDfU32
Tagk4j1L8tR67ctqDLSo49ZVCjCi2JCdLCAIjiE7k/47u2GqIMCiNrvlRmoY6uTfL/85ARvVFV7P
AG+zJeclbqaQMoRqGSIBGdYdwtWB1hQYdLXuS1KaznjcSwTX7Wy6P9QjzrLhcoLqYWVW9xUviM/7
QB88wPAeNBqaBeBW2H5ziKKt5uJWycQFz48KQYjKY3Y1x4K3If5u2WqiTksFl/RjVhFDK1UwXb5F
TEdqqo2hhba0U2LqGQ+u9+d4Rn3x48rEV6jB5/qC5udISz3KvsaqUU4bvGfklFdBX/ok4sZ7x+cH
SqYee4Tz5HYT2Eh4NIvQaBgSHvj4TJ2StoO3ClAenn4s34o52Fga0rHBj354qW1/0AxbLfI7Tux8
beY/RPkWt6bTOwVwzZNFy863E7xgpkEqECyI0XsYJIAUYFucvC0wSA8IBf2/izy7mhKkMHRnzAmK
Sn1TwOjV7PVpggm2A2YNCgT8Pcnds7I9bbWIQQub3kHgQfa+ZeaE/6ZjhIDbg+UMoQzHdbFS+8kL
d8bNyDBrVtqGNBbGHfkNsiYRnpa6dvXNozD/YiqkJUYadeQ27WLIAt1fkclJrzZCY6j0llq0we9i
3tnNl60a5qznndkUuAG+IVGC/vv+a58ygbjEEmFSER3zvcj0lWcIcxmQcWqqMherpgU9PQYAkaDq
xzfWsaXdOJOfGHlUvgxRXNDJVetk/uVGkgb7hm6EfHqEVzSmugeI02TmkOuFVQn31HhQhQqrty0y
0ENX/6dySqYXrUQt1GoerYa5CJVZwZP9uikEpA/tccdDnRrFTfPbmpHbdMS9zKrT6nnQLZPg13Ou
cU09aE2+CdK7hrvjbgMZKojgVnNX/+guznMCZnK/V+7khoadL+PCqRyOl7FJaWzhzG4Yda0g15XO
+0hlF0CYrfvhFBg30vSwHzepxKhrpDyWmYAOGcZ2DxTQzKv7ahqi6Tw8i2scBTsMTiWiBjjyaSEu
QuhXxy6YfCofE5sWnZmblEYeaYjF7JNlzYaMvY/j3XtDs9YAe3ByIrcUS6oh6Acxmoa3GixxWElU
abWGtn0N98Nx07eM+qFwtF0b4UV7F10tsXdivh50LPR/+GF6M+GuMBsQm3ONKQLGNOuYT96OZ0QO
Owek/ybZc6Vd3Ib1Jrg+G1WSaJ0bGEwp0xrQ6eEaonhHQLTyP+YRX3YoV3kvpwZ1e8BxU0H3KTMF
I/g8LSgUa2hL5Fh9wHoWLhIoLSqDRwXVA8TTQkrvk1+slB60Nuv0mooR6X9mdCCb8y/zEsN5Zrn1
4XodHMDdl0s4ibKBzwXqS3xRrfbVbqenul7iu795LE8yHGMtkgIIIcd+S/5VuDcphvSNC5faAOoi
tfQaXnOF9mNpzd/R/5mM95bc09kX/Zib5jhXQxX1uBPk3+9LDEGhkWqJ/A3104RlO48gyMYDLfbS
Cf3xZuQYYJ9+UELVSSPK57duNrSPwgFQSMhJgBgCjHIKWtCOYRVKTsRY6w/0ALvXLlqwbUxwUZxd
xlnRs643S7AAdZGNW5gRP3aiRKlopSlGH5mG+utr2mk+5ZDj8+/zSk9WMvuTp6ZycljzZlWxYbDv
BJsqsOMKVT2bXHRP2RKbmX4U9o5vX3aJiHelt1mfiXc5+c5Sfop/7CcKZK59bheq9iOmfzfHb4QD
A+nL76POki7YIrCl1aLw9hj2GcYDrXkhjqRKGYpoqCMwOgpqWNVANReY5arHgRcZkoYtVSwisFEr
pxIgm9Fj3p3xq6ZttuavkiKjHD2JDtCPlIwmUha6yzPh6XkL6HDxpu4W7gynmQvgGTG1vcHnWyjD
JA/JRcYRvXnVhn3eFzwKq6Br46gzgoohFMHJYDu0ZYwzp/8+ZvpA8o8LXvZeWXE5oMoYwyrNdhiZ
9GfGHZucoMFQ0xoErvlQOLdkVW6dheDADtGp+knDzbuNZZZIzk4GfpmNu5nGh5VyfycIiNN2LuPB
UKGEJScIwA9tJg/3hnXJnkZgL6bc5DkhIbJdneZZGIz+XSUSc44Tc2oY3C0lTqgvmyLCUNJkYUNY
dpFf81byelZhWlnnT9vmFVOIvUUNyGUuLusVsH8iTOAJKIzHpuvErDqcXMF7TEgtjURkIuq4FzdI
dUdTwYTf6P6e9XO1rpbnaLTAX7I4HQyDKoG42hKfLfLW0R5EjVGgVXFwwcgPk/OikDazOhGv+EqM
xAK3Uy4yXbriSKlZ/SI74E1Q+1BmbfNq1eoUZlEjwZmyhKB3rqcy4cr/BahUtSylycVBrcBpTL0X
w0UHYQPmuLqW9OQ3aPTyCDC/I/nhCAs74+Nlnfwd1GCb3SB26qNHXu1w0DE04HMMxRS0FeblZx0F
7FxaRujke+dbxPgNrZKrHuj3qc+wb3dzKtbuneXa6d7UEvowL0LfYC9Cf6TVZJKNckW5qPHStPsY
X9CjqXC4LH0yihZt0vEsV3LcLfaO7C3cFKUFqnyRtyKqPeOxGE5m1ODuJqo/vMLpymZLHhgwH+6d
eVIbTrkseq7G6o1PkSvmeD8p324fDB2/iTEJjjhVwbzbVZV+c8ndt74F8FudUQZFlZN1SEKlnjZJ
hTGaN/+cpOwgLQAHqbbegBsUIWxAsvL6uzHsR2io/QFR7+hVy0Pjs7Ls5qq71yHDu/dZV+c3SHcu
8Cm0eIjPi8NYhwZ2S8F/0iwseFSTkojEePyjkVcvndbnhUj/ONJawZF75dVvPzFEP2Ob/XyzfR51
zlPUgi04zQyzZ4F6h7gcZDm/X4+tJRPov8HeSkI+fAhSM2cl6lcLo0AV8Z3FFQWaQmKin2MJIEAW
5L1IvI+Vt9eCBqYJcGMh+0192swXPAOhDdjoYw86fwIFo4z0ihvG1R20vyy9PrgYwjUkojtAdpur
Xj/taF9/wsjEsPHp87hSkrnp/AJYfD6M6hQwe6dYouDE7rwGMgfqR9jyo+16KcgCCImgRbFeoHs2
XdFCQnIU1LIM6QdgcmUCWeCoVevdPY0tu3yMQ/FXcJDtf58mNoHQIxmAv8VIBiazQedlBOhiZjEF
PGICv69OGmS4MMVxOfHU6R5tqLmughzxUFR4rDmvL5Iyj5/fDOnWs1FCD37lkk2CSp4VopeE+r61
hhA4O04URCYHIVg6tgswBm61xI/gyOHIKxl+sZ/X6XNdsHnbv9PlGPly38zPqffVkUKfkNLGC6V3
rlpawYwhhaicsE1beQ3MlQqu6aVxLj1F+kDE7HvGcUB/x8XrQRyEpnKR1+iqRnHVr1X603uczQCq
8fOyTrhATEPkvh8BM6STXjX9Oej3/FXlj0j+2/lxLRe7BFVDNPeNJ73CqdjcNvfiDZGT0GDZyQuK
pbW42AlcB0kJkfFYcXjXtPNN4FtgtftTxtqhE+f9UOUFFvNMq5+9/Y/vHI0faXYxeANzSszuYwiJ
cbd6ULbfUOQldaJiaEanaNT5VtLRLKthJ0ymmv1qF4RntXZvvhKebkYS9S4/cCEkqh4iv1nduKt+
qpOlM6vsxGyXhTcmNa2hKaeBsWh1UpT1ALJQ/FaJWQSjyb8593zICMrJFLhxrBveBQNwBecYZrSj
78j1wnJEpNWaRMR7+sAVJ2TSDOrjN5TLNg+qREio8rFCn4T3HuTTINN84NOFpggf2CLyf3CYEblX
JDyY7NdLs2RBlsWnzv5TkMCMRGIGBVJGGiEdgdMFcZUn1UFwRbN7oc1SOhQi8dg5qWYMUtvNZlDX
8M6buk2zg09e2PeEAuWi1ZsuultIeQScl3e01ZJnb7j/WnSnUIwNOmTlg4qyjEHqfkvbvyEkbVoV
NrJ8NKxAffyXHM/iZBibUFj0PSXUF+c1ryJe1MQhCZtww/IDvlw+18b4L5lUclgW7rsBxm+cUcZN
NInp92Zdbt/d296T0xq4kLSeM+mag/PXcbAofAIxw7YbobTbsYxl3jjFF55oYf0YBhgP0lEuFSgt
xPFNXRMCsIA/SBN0p6pvIuRQR09smnns9xcU+U7dYE3FvnQZSYSeMv+TCo9f2iDV9QXn7bsqZjiw
5AWZx74iYZ7I/qOfWP4q7BHCmZdLd5c89kvh8wbNOcLi2799QTf1CnjrAZMNHKwUfFhjwfRRocUY
4oaQa2PRRcyRDMX9Lfii0lx+4oHMsxt/64/cz5vZs+4rqlKX2xSeeON8up4SSDWpX7TP4Nit4PnW
KsLn+6yeQyViiC5OkkEMiJs88bD0idaRhI9iNmW2jAdo9kSXGcNVWA1TCm1zIMpyfZDhKTij9Qv+
dpdtUT/XjrN/o1mXujGFb2XHgaJsJ0PGHOpRaRraggtcAZE/3vybpuijyDJvv5KXvmFtsa8pu7HP
ndSwRlDTLOrmq1IFtRF21SRttnc2bgmuzfOHSHsPn6LqcTQSw+uxBLEFhwkaEbXDU7uWhCkC+RYc
YPKcPrXwRZEi675PHlpG2Cujw1XhrI7ZS8oTGoQOQLAiCAXHGBuAI9jJtwa32jQQUvNKEvQP9+hH
A27zph5YTOD3cY4LaAi5Yb6SpPAHEqMBalkPnrCGWf10fO+xRpdqhmPDqtXWVL4bxCqBCDUTFfH1
fflxTmwj2xED29BanB79VYBchLhht74lBiLiGaYBdUB04sZSNhCNAeyMCBKhCqXeIcxfZ9bV/Div
03JTN+dNxorBkx+NxhopHjkf/uMXdpEZDsCiy93trfY3EkE9rYAZ7UrO0nm8QFBWDRGkxBPVsFyu
w4M/RZIzXVijNnIjYwZpIZ2jtaOw5wPEY26VXBJMiJnVcm+9mx6RsaLRKxz40AYlv61IEd9wYxU3
mJ53YyLrTfc9VUWbtqVBykUvkApiB/T77TPM6PZXzPp3MTR6lssEU7xMI3uEwiS+VHMPf+/ofWD1
ICEMCeYE5wHxx+t9Rd3nL0Qp9ss3jkWEBWRpnEAWZrlsFgl8PPRysJveZAA1OusJdxd6WkqJS1Iz
fmgw+MvpafGda4hjnTutvDBqKojUfhL31rOFZC3SAWKA2rV16TruRpJTKoVIb2BFofpuyhFZr3Sw
04RgT39U2Or1tSZh5HsjD+UXq2961oshjMkuXNKv0faUZD4CtHwTqTiVMTsxDue5QrkQDS9TfrHX
ea1dhcIfqOa2NwAOzfl7wKUyyXXqTaN3OMknRKCFNmKUd4O8ovaAYrYyyKqK/Haeg2Ck8djFEqKG
7TdIi/1xA0E1AbQqKdw41RFX9mDql3YTkgvAGsnIAV12XEJMZDNdpEAAQYD5DnbAx/P/Myqi/o+/
+tpYIZWoUH1Nm7vIFLaP87RtFHtsR4Nj4Y40K8BQZ2EN1Zc3sGGytuGyR3HyyttcF7iP4gXYD0kv
8QTxYYxLooGpsfDw7GJMiVKbemRbV0uhYPFG1MyDJPKdVeI1QJ77TJ5TENAey8q4ua0secBhx4Tv
KZf6NCa+qya7vcIcbNpxTgya+n+q51Do5V+f+ltGD06DvzVPPoOy3BhqnYbQ632+wZE6clZkZSXT
/Q3CeoDnYyMLY1XE8cE//lIiCq2yGZjqnWeHcMqy731QzJyPNofFdKQ/uxqKIjXpznKS2NAPdyp4
8HNH/S+g+46Vp+LVUKY5caQY+bIhEbXIYHnWoZhNdvyhaq2ICaIEa2t+7VJ2iIJGcLTKEexEgg72
UvTrB/ngZdViEUQGdMZLfQ17CkLnh03Yx5sh0XOexYUwZPYK1BtyV7qoC/VZKq1uw6zLKnLdrub7
q524pXTXrGKqxyF5Mn4RIynjbmn7UR8YY55/8o1lWEkS/WheLUxYAKCvuzp7M2qpv3opkgWhT222
3zDQhiSfEwnwY/+rM+0c/DwNs+bwrSHmpulxtkf8vYwOGNXldDGjXOiz/+0TUZfQhIzA/7yFV+Hl
0u6WAoXng1OFS9AxmdHztw6DREy0w8200kGTHBEXv8asSZic+IpWkHR/fvoDnvO887N00wuEjV+d
81ria+WogL6V+TT6KBjujVCBudh6ZbndOpt2Mo5jCbm4magAPpjL3knMFNxfCb/oFlsXUEkJvqiL
97DnfW83VVnKkcTuq78IDJRwWchGcCqfnerVG9SYa/dPZbOQmNU4kH6k1wi+w35MTYVTRzyx6CKO
C/jDo4I7pGI1Xk/fhNduyMxXqhnGqdTjlfd4rkQmThNIhELRx6B2e5p8aZVskr68wX3o/yEaQDs7
FEApyMxF4cVOKzqvY3QZ8xAAx+aN3XqOybZYYqkGnffm80y6gPksDlXIi9e0PLKn8NSwFmx/lsHe
Q0HRgtNf1NMiZs6YP4ip7LBKpHK4j0doVVTTp0AW61bP/ri9sDiN0aYFR97yXY92yAoqCvgf1NFH
gjF/PkKMsdunzzfFYwgrsS8KcXfoWhUg1osJAoSdJdtxvm/qkPte/mwLpjhQl3TdWfvDxcz8MIA8
lrGhBHw2XeosewpG/pbLZN13cDSl4y9lFarrbyp24W7Nt7/GQO7vGJDsJVzfdK/3tu1VXu/6c8cf
gRCDjG9hXOVCHBb04VFtGYi6kJgqCP2+HvEyGhy9s8hKmu5DPKDI9WCaSj/MrqnJyykkIscgqlis
H52qTdAz8fFIa2q/vvTe68FJ1mYzSzenQ0cOvQ2TwCpLshSynlPWE9LI4ZzpFKXgT8+zD3z+YfzC
eJ4TOEn8/F4WX/rEz1Q3ComvCS/nR9vTQGJzVifxDgU9ZZ/hwbXOCfIugFedvs7CyWabyBrq6NqE
EJQbLT2QHS8TJaDheJcfsXrGWYxCnhh7Cnz4kTrm5/vEIg6ZtFwTwy50yNrPsQo14WKBUnK0cxPN
JTPfCRbh18rm2K55UJqLmrQxOgyywszexUtdU98B/B8BU7eACUi3HvOwTgOr5qSDnF0HYoprnK5s
ZHHf2Cx+UUeFZSiSySGxpSWpysZQl1zNku+VaPsojYaVgqA/8/8ILNla+SD0DFDl3U8uPc2+IUkA
+1SqhDPpTPFnKeO6dmQgOD8ToHDzkAJn/xKVgMuT+k93/pweGyU2sb0VZubGXS//xblg82OEsynp
0i6FkrSiVuSM/M6VLQINnP/YFszVpyNpRWNGkUcfNkTkqkvwl4CHOMtFTa2aSbtqedImkbIASF1E
MFr9HyZtJ8oK8MzX5NSbVthnnKHKcZLQd84ulJVtYhVeiPvjp/q1c2PPmpEhLwhHk1KgZYq4JqrD
9rjB/T+h54rzlziQ3vb60pLe+O7b2sVbpai2sXDm1BFFafMgMaORZljqAwxUHZzs2+STLsvlq8aH
+heu+Tk8jgJFb0kYIiMCbOwP81/RytijwO8NT1QpCBNAwWHRAQnKzx943pNxSPcZoLWXHcVAzzpZ
YpQ3x0fWHkpJXeUPtDGCn4gVhEirUd8upIDH5u3BJlXnsytZ4mKtVJIoxre+3peNSagrazRE3dhs
ytsTYSVnOFevaE1ZUKuK7gf9jAg+lydudgoTiM+hWH9lKdd2VUiNPhCNFx9gJhIiicrie7Ht+QmZ
rFgZfJZ5FibH6eLWjtpsWC2d5bWbYBJauRKvOWh0E6TxgziEVzmczBbtrdg3Ep+E/SGUSsT8Azbp
RlSKThLfg1+3IaNUonlSv2L7hkCCHz4gnLeeJSo96VeWy3PQIaPiLyzXy8BLTQlxqfn9cg/jOFu1
OmTq7bzbBmWDFRktdhJFRMU48RIuY5j77wRMv58tEFuV7OT1NvNP09BJIFpanSjf81lyGy7LDbqc
mXUWe8tCvSfg/lXSK+dHYjGj4VTW3wbWlwvIee9kuI+p/nmc1c1L5oc5jM+oR8CBbHSOXHRnMFZu
PRp3ROY1pyX4ypiUtj6NJR4ru5dYexr/5rNKKVaX4Xl94/SjEwTBiANcmNPSG74g84JPcuFVjDxs
+vkJuz+ZU1hgciAi3pH7m+QW51t+fn6dBBPNCoe39FDNDaIlC+CZWMB2qoVvRr9mntX2U97+p4QI
roNmpFRnrHe0967Kok8e0D/0XeGPKxXMZjyvuCnVw4Wb32Q9ydd2Oe7RGlcAKpZ69tXuST2A+Kjb
K4QpKmX85PwCEpnS3DJqlUBhZx/EkUwYXjGvDNhhpzRW0mHtnuoTw15CPBYI5Pt60Yumrlli/2AX
2+9jFxbK3oh2NZ9+iI6Lna62TT/TPSpBOkcLxMkvfj9EYbCXtTLLcQcbYIIpkGuAOzV3Yqk2+W9X
wuA0YgEm6Oz4dMClDolrZ72Cdu/Hk3H9/NAYmabTx1WfYZSQsyK6kdoUkjvTJ0F4HnIM7C/oM0c1
QGyCNWe6MW1/3mLDwwEDLeFjvH8ll/ta3CwPbyJWmsFSQKQsPFDa5ZPysYe0ftZ/kghwkaZ4i8N5
5DsoywLlbvlXhLfz7CGwhCrGmkaMQPaV3Kq4VHmLEbUQfhIoNeprYxRlVKaRNdlcNXHh5DptDeRs
usvq8LiyvJ2quaVVkdx6Or7B3fJjJn6ePHl2M/4a6rEL7IqOXEMMkTvzNiqcEb9aQQygZTfXZARp
k2wQUdWFlH3tqJ0brhdUyPPxE/XTlEv4RRzvxgFjFie26nSIGRL4ONhR/tGDqiaiqykJ/GKSQOhX
DuD8Wr7DYTiP3T8CnKpTWvMOrMngvdQiyuhM+v1WybBTQcG63b/mxpe5slW/g8Ez0hfqjQcEjBfV
tI+NEOA3Yysp97WdUJB0blhfSbRXUzGNNhZ7pcFrmfm39XU33QgmVBaeiDTTRm1jVB2/99ywwVXX
Hmny62gN5JUqbeO+nNb16hXnxamnIdsaMUC5S11tPcrpOuvyYtwJU4rkxrYCXYPAB0HKqfbZX9oB
k9+5wwBckgBbvuPRDBuKBXI3KS6QDdMCn1Su4zsSG1IOa2BqGn10pSQkJZV/+LDQ0TLwAbdjk77F
06KDbsOzFZd8H5imxO+hr4lcttYZUCWtYTMh1+zM+j/gcXsQ2U5T7/NtTTxE23LdnYSGsbVcy+i1
9r0Df9YS9SdSEpPQLPAuxE2HKc+N0hp8ebrvgcspxo3yt/XRA+RourIUn7yXRTrzxsrBLGpxzIhk
8Mb/7e61gdK421kK5L+BbB5dCX5lYYtHXwaGOuorislHGBEjEtJq6jmSWLabnXgXECOBhsKGw8hp
ccs86Zqfc+uKntVWTos1W7VBgY9R/BLhtLOpgfRZCIofvwqvKXrONGVbKrKIRhQSMiToZ+OOfOX5
rRXBa9BewXI72WBPBNZFe7WXlzGe6R9Swbz7+ilfBJjkwYa02k34yA78fVeag5xbLyYJcqW0ySMq
NqZ9nu3g3pC+26vpOxo+nHeAujdK9Hcny226Z/3jjmaIxTkLOB8nbaB7Ad2c2UGf1LmkxvMEs7PV
9o195ptAlu21z3oxqrBI/pYUysOMBBHvxEZ8ZHyjg2NWuzwsYDsVGwYSWLK2EOUY/EaNYX9St5H1
T/e/jGNJe0u5Nx1ZvPoBrJAgTIUH5TYTxsSYwvT9fhqQCEGa6xpKNcyiS8ZM0HhksJB0X+5sPS1X
b8mBuTPOE9hpDde86UCgl3STwvLbK9+yiF4czNTeXLUin4vNSXYuQVjkE5oxc0RCYJqLjHe91lH6
WqMIldbVDtb6qEpIC5jDDcGMPQmBsxdsromN9btDw+/WavHGnuqBaq7f+dD6iHlSIaS1RpMB/eJP
kIUqXa7mHdxRH6BBEYeqD5sQs3znbu0lKzjuQ9GNlF3mNTuKK5cFj2Zy0kOEFoHR2X5QCUMwgrwV
gw1n/481PQld3s0XCDguxDhMc/hiWHi0GQk0BxOCJeO4PJRkcx/9jz5G/n1LJ/gOYaZVI+l+WPzs
lIKp3S94Lu9+3dc0vEmaJVkPooE4Y8e4NixY339INGUqtmXMRuAYWGpikBca23ySxsORLvTvbaG4
3aAwosaZOHtSswRPPp7MUcb27JHuZPxvj7OxewyQsz8GGhqvc5PS0eFn40VDkChNvX7R8cDWnlQH
SFmbF62Vu+d1MhMniYEVcxWSIDtW9s++Je4yjSAulQsgGtYFmfRq2p5/n3MBlEbMayAsDyZrQesp
lLGtmy+LxMEXpn+/uxV9e1d3pn6UjgCYNOq4Qeo8qv4RPQ+ohk9TQeeCdL4fNgxoVeefmuXNnrau
kxswthcIeHHBn0mfQZrGabqUPHJI7VaQc3mzrxioeV7+sgZWJRj1ZtH7ouqa2Gx/bYFfcM/1dkgf
a4iaLwKFIQRe6joonDwowg9WPF3x+Tdw6WxYJIpdTC/IrrSgjVWPuC0qkoPdGUXcLeOKLyK2tl3R
MLWqBvkEN0ERgu5ncVzzM/xgErZXi/FG6i/PX15byOVa7QR4ezLBf88UL/USSKnYL3wEgCn38rmL
frkmLVyatE0PJeJatqRMTQcX3CXzgZ+uR9l1UqBGkS3NIzHKQf15XRl95xWaFKPQbFI8vjAEO+4M
JQjeE6Gemra6rQSrOLqdl9TerMTmLDMjcqZ1P6d+dXoLw8e59ADmRlzBlDgRSedtt/lqS/tKFT5P
WWueTMQgYtlqMDVVYoS2xHP2ZF2MWfC0rnCAXA6dq2Vi5nfEOPW+RzIt8h5YnVayRJ5R/tGonUS2
yyR7wSfGfYnYqOzxrtE00vZuz2bdyKYC+XtHuaCE57VvOhdnPBCOIRcxeNlHBmjQugOoxiCbc6Km
REyZgDzwW3lpuX+EgWDdKeY1YQWG51pXELGgNziblDcEyCWsyPUJ5r9ygn0DnALyWjD03K/6AQQh
63YNKA/1P64isNYxyMuVB5Qy/hBGIuX1iTIkEpgCXuy9enQX83CQ/1uXvJ9mV2RwhtHrxd2h75rE
C980UUMQDXs2eOjb6vdmxWgFlMAfJmkGj9jk8swOQs7VqhgNJIRqL0dY39TZo1nz5YSS6SSVrgOu
PZQRZNiLjt4WvpTl2pOFWUg2ZNB95D+Io/oVs8rLAszO6KtrkEmlkqiHbSPGwdcHCjbGmxR32aNw
hj+U44u5IZNcHn9VBf7oIc1HG9chRCuPupOy2x8zhWZga7P9xQ4JGz+N5Fcf7fG/74YgBoOGfG1z
JXGQXcKJwK7Q4UjCbesYGrn+U8BVTvMsKjUC5I7VGGp6mac5b5ztoeWXF9z6fldUixrurxBJogGq
bL9woL3/74W80m7OZEVxnYWSRtQWGPGyoLuzyvA8h2afo4Mgr6TlyIGfTzRwScA7nqLJH7c3otwh
mlryYIp9iHU7XMy++19ppC+GzA9RAKepsq8ONVapjB5Te3NA8EiVltX6IhPkwGrkGNMnd7syK12g
R/1Q0fNLnJugzSZCRg7IFEmIQab6S2Fcc2gley08uz7Tv7D0RLG9Xr4rrWe6l0vsZYUEIYGbKogj
HcAMdaRYqhZYgwHd6lrYxNy41DbNR/fLSZzhRzFo0rugZ7Xb8NIMG111vJdl1Tm7LBz+iZCwXeiO
CPWOglcp/0+4uARQOXFe/pITbSYPWqFUotCYAc5WstdLw3ZhdaYbvIsuY1dJ/kiwo5QwHZtloTDN
Q4g6sp6p1L4imKo3gNtj22Ifp/Xiont6RxUV9TLoh5l3+IrdXKvETIpTJzv+o+aLE+QhOZNY357F
xmzEZiuur1ipOFAG9oImMyArMFZtB4rTLTE0HPFK5iBYmufTHTEcYIceWPWRpOhLq3ieFQAEZ65I
Bmbx7Zh7MdNxAdF4V9kKJLVrOZmVheH0/gltEhSZqiKNk7qWUbtlruUa3NaG+npc1Gm3jQG0brPp
TXd5/T3Q1UKDLzk47291i2v2oSgYSQkYjV6V1mXZllNpdIR9JZMsgIPkcJcuWx5CbZyVwjl+3pGO
9x0xdXe8V2x6P2g7ZCtK98ZSyy4I12N/I77DapXCw26XFRbzBui3utRYBwAXp3+RC55+VSPFCiew
7o8HxaSzKo7TIQGW93UHktKVuVOQ4oPGMK1XyZ0jmc0HtT/uLkKiUjPz+0rzBVT9xvDBRY9uvFmM
YWf7SWxY8kU0xRieXflVtM5V2X+wHjqGbG30vzyz8LACeWhN9tmOY0++qIcEwpbg94+MQs3/86Se
/pX8gMtd66KtWsdLEoJ8c67Eho972jgjsJ6WvhP/Iu77sf4B8as31DDDAEZIrfEeXB5xm2csBx7e
/ZZobzz1whxM3JSrg1brFlLISTCXZu0JXGZ6SkNJbvgUxfim40MNMjRRItfqwr8wnWi/4hMbkRFY
RZOaR4W04PA2R5sUVmBxfoAm0j4+XrmAPh3tRXcvdaTgQ/1F45HtBNaGlTvdlJZsQwTstsOPtd+B
Qe6IwO0NAHKwPiUxKPX7o/r/J4NKYp8wyRM5m3v8NSilz93sCvEVzK6dl2ZYpN4E2LO4oKLdfyPH
R2olXRCFQI8HdAur//c7HOgiDbF9iWUVpB5Fny7OckTxXKmrvZLvTD5xdmIasISdtXE6SKK8YOJR
RqOSZKrEV4eN0yTKA3EMs14iWMPPvUbpXcfuaIFS2ZybNrz5JVjRwyyThS6gAy1UQp71fC57g8pz
x5aQEpmnquTevHUGqS/xUMyg2hMsROl9AAMHZHOs2vCb+wzEwuOyxqfPL7t8z2lXoJ4JMfY6/Bwi
OxFcrdjiP2FF1hSivAhn7POaaNK71DQzpxa7GqD0p5/+fMXikn+q3ZnIcTXl13KBd9iNBn3yuDWr
ZusDQuz1J8qCo+pElPWWD84JLj6XgFbyH0lFIncNweo2n+7rNBwfOhMVckEgBU6l+sUeGOlc+y9d
yKOFU0tlHI/8425m991IiTaEX4TrUIGuBylmT0kVyikGWhEFSQdnCwC0lM/3WORmYYzCe3tKXxtk
xHpDt6ug8ctKjXFYxTH/3nhM5fXtii+s3g1L24S9vUaHuUjrTlx/MZlJPyM5AYAT16nxnm3TueAf
rqhUtNrvue55Mu3MxvczwBe//1QRxmi69Vfd7J+vqf7gWO2TU3RHeYIC7TSsTLZsG1YMEpZoEWn1
9xqViqEjxOMeZXn2UKucxxObieXX3Zrj+2tP/uo9MASDTNpV2Qiyl0Uj50a+pXBySg+HsJrJ4skj
5JpAjgEN0pazLFLikkh5ZcU2SVuXXRWI+MtwafEYJLfTrhpI9zCz6sS6U/o654E67X9FRUV47m4e
Vt/SnJlE8Y6TD5dCuAz1fyuqIp07XuXXYH1x7pV8TSO3FHsNMysEz8s0jiNaQiKSHq7TwbqeBHuM
UGS5+OVNawurEwJRE8G73dLJ0zMrehnR+cJC1d2k5/77PWmXAKK0dBs2MmTWW2zoGSqlzMY+4KHD
brkviHp+g047jul0+AwNIaXsT8C6M5CMBs0XAaEB0PiqRGqYuQEZSxlzWI9JqRRerxWJVzpPVo8e
zZpJ4ZMo0PE3KYQyAV2x+d2vUU3h3kaBrNth9pbzBYEGp/Ia58WuYKxdOEjNqbuqD/11GgboKxkL
yujZNyaW2wAsllmSt/WYmzTVhvl5Hm76OyLmQ6VIB9uKe8gZQ5uavJfLxgac15jB5WbE09juBtMq
xu0E1Bc3Orss37C3JyctkiQld+kwwT4Y8z5oSeCnSzMxwCg7cmtzRPkPFRbYwB6yd1nSercmRqOj
9RDlcxtQkBqt1zrmj9Lu6m3v9VjjlhYJNwBZvjN+fbNpOR89wXkBhH4HRiCVcWhinyxen6b6SmI0
DZfmfAP1hNOJe76iu0JtOzNK4oOjARKqt/P7cvRTQszydCVj+Z5Bb+/XKFoOBipeeCAxNvRPA2ZE
oEjfbBOmSjKRctfsRKnXzYE6EtLiOfS8NLTKVNrVGUkpmnH8VWxoLuvyq4ksYyIMWzLVnUsV+AR3
TUrLInIeSMeuUQxb6iM3M3xEy1yFLNst69U+dgsjWhTzxeAzqhWqq7182SEZXKaYyzoOI2CeavSX
hoq7ux7a9z7N3upZ/5MqIeVfJj7yECaAZowkCmD7teVNRn+zEPdgBZmJLRG5unY/YQuyDJiwIRYc
ACdTb4sYRPeJlX1PEz57dtlhiPkRsoa+yaUnzJquzAXwn/QbT8yDnFF19zdIkERTfAB8WHfFCe5w
5LNAVFWdpKRtqGEdJr+26e94cad8C+EPrZqZLTJ268f7lfDdHeqsOwxf4XUj6xgzZpXUEt1zHldi
8vM9scODRI3GqJSymqk7ZeudFh5VUwH2Z79yc1rzE3VjzMnxEmbrecChCL0hVYrecRaGzO8r6/wC
IhczQCmGbZNIA9XMnUmjeXwvgAXBm62UVXcDyChj41bMKUqMuzc7vVaNs8yzU2h6INWxjHwhbMuv
E3f8sqey3PLFWnRSIfz4Mx1cIviPezNVE8+zJEKRE1tgby7YCOEln7S/WMk8+NA9XEk0hfaKNmLb
qIC52gsBorSFzwIwKcD6sJwPdITgIrYEEzcHRHkGxZkULhcIX8oDXexpcciGfUocYZF/tgD8bgVr
nmgu2wAW0hDl5UNLU0uRCbMrvmEcJqnb8MYVg0Ula+zFAKLkriDprze1k+E3Fad8PsUT5y9xtxUA
JgZHItWI4moyZzytAhoeY0wV0x5dEuJh+ipPA4F3umS393LbGdNBvEo4yH7sw0H0gZhlyLH0UUqx
qibREcAcU1dJHnlUMrk4I0xPQ9tCwUAfo5mnhL8uJgfPF4R79fMgZSwGKpczPqz4pXw4AJD20qDw
VAYF0UEejaxNPLz+Sriny7Pt2Vifz5iAv/Zm0WvzPYO1d2T4cMm6XZ8RqHxna0vaeqJIlT+C1vdn
Bcdn03ypp19gKUnsGzPsLTMqk/s3m6+iGObsJmM8ze8XnMjvMTlxf27SkODmvb7SQaiCcaAWDIxR
PkAbxMwNzRATw31KARzGcBcQHx8h+oNNh8tW4SngytEpnKEmvHFH+Z92k82X/HPi/STkgvjXqZk3
0BIyW4VdFjv+byu5vjJ3z8wocvzVDm8MXhu5DNz6OgWK9YSq6HvvGgPVPDxrKAMn+ESXamDu+fWs
Kuvr67GiNsu2LBdTOWY1qkH94fmBVNpFd2Xho02A9PIgVE73rr2yPLy2DbuZNEjtLjtDX21v53Cx
bv/AGxHVnSPiRRHnYxN63Fs6aOMoihhUiyg/FmYLsBrPTAd7gbu/V7qYJZxtcqqFFMqih75EChwx
R2vWuYCa1wnGfRe9e3Lh5YN6EIGgiaqpmUm1DuMCY79MLrx0niVxP3mYt1ayaH0VimAvZOvCv8WT
GAZPOA+oSOPFgDVa40ryD1k9+M2oKBI9wLvytDLqbesT0/IaZjexBFt6msKIP2mJVi1AS/oR8Cko
soiS3lBDmGG5lvfAaZx9ekZkimgyKJzxEJGAcRmR6UR4swe3YeFfeJZBQQBKVttftL5LjF4F+tBJ
BBX5FhXRDBOOTHn1QyqZLd9LiG12KNKjN2PjiFdsuNYh//BkBhJkKfZ63IJ9MZGKNCUbR3J4XEYM
nmC1i8D/v6R2fdFE8XRjQ3v+ixfh1cIejgY+w486sDYNl/RyHR5lTN2icA/yzjrht+koXkf/iJc6
jpZ+TSL7tGS/r+VCRFi3UqCgWdoGntkFlXMPh3nTzFLkFSW+pVstjW1tA6SF2BUiZW4UcvgyQuur
9Xzd/Al7f9YQgwXVqP51EG/BeX9NrSCEn9R2/2OlR0PyqtAyIt9B83j62KvvexAWwfpCsxHCpEsc
GLNw1GW4M0DlDILiORS4upI2YA1DAWme6lBpnLHKlXMjEk7PmN4MTAcgRqJ6FN9NUxV4JEcV0WMV
5b2E0otDoHZiGjnqB6Sa+0IVv87jg/Ge0xfMkGo1JCE9VbN6qME/iLEfzj0cBeBeY0vOgXedqoqG
gwpSiVmsrbi2Xa+phiI4mVC8gY8kz0bI9VZ6tap6hoUCKPzVZ4JR3BSB24E7Sic/vnYdsqHQVsRi
KazqMMtjwXQGIJLpVzqUCh0nF3sr5zK7dsB4245O6XxvTALS4VGYJVHunA8ZcisQhNUpul1bZEGR
wfZQ/39QYCBAiJG04RxfCTtuUO6tGeh4tw1v+3odrQmNp5KeiD6GcfIIDzxos7qYNqd3bxR0tI7I
oA6/qBvpDJCbsx6A182EMlGvs6nbhP9kp8xPurUZ0fJTWt3jSQNhbdnMMFwUO3Un3kAtStyaNi/a
lpGDim4xGcPKlIMHr8aDdmieKuXdlEEgVNR8gv5yzVAtziCaBk2HFRE0qAsPNSOAg1yfqauo8gbu
CfrttzN8v+dNtT6xTVxXTmPS+816fLi3FwVMct2/2usOEoTJAyfLb0aAw4J7Jr8srA7Pzhcb5HhP
EicSfMhoZ/B+SrDoqyBeOD7WClS8V7089KIzKeEFqDf3zWL9mrTt/gl7JnIP2/9THCn8yWyn4iQG
d8xIN3jqoT/4fWUQSeZ2MVgY6Yshfy/13GI57vT+jALJFCS0OtAJzD1TdTVxOYdglPbHDais7ibZ
A7uhxJbsWvLBi/CI04J1QkmBLMGbqEGX8AN5Bl1MBl+vC8PvDEoF3HEwIbV7w0wlTSxAMnXVfQ2L
rZcPpRvayDjJx+Cam7mLIhOhQauGXIQPkiVoeyQ0I5fsWGD/MYelvaLdImB6gjxOG65+ox76bHXz
D991RRg8QvsVeOhjYudfI2Ze1bM/T1INZE0gUxMtwNhfrqnTrMBpQcQywMUbHfzVn8cmjKCjIYIC
LQzju2Uk8+subEcj1zdVYZYt3i+FYHcJ5qBSDVkcpuVGrZ9/vrW8DoAJ9DdVVG0INvQSVeQ1DZHz
CEncbP6TioIj6GMi8P48qdRhMzf+Ys7mZzzWq7HcdI7Ui3Zlg8sqfG9gwz5vNET1uOOgTeTvN7nM
dA3Kc+pY+PkPcgb9psGM/n24XddzXBHgKwQtIm2lJurwgAHRhK+Fvpr7akhxtzWfZ+GHM41gTk8q
SlIb6f/uVCKovOdvP4EmlskbbUAPqLrwBg9LphyerMUZ1i++Gvcpyz4Yq6m9igD/0NZe/rlk564C
cFCC/q2doNwo1MMjtEFDvHI5cGu5vK7+eziRiAbPBvepSBI+q2b3s4fRu6+79iySAhV95Z5suYLg
ZgqylTosAnhfwbExrdL3CJvr0ocZCo7mAS5Ikq1Vi7Tb0469GagIFMkeWUr2tMGUIlcFHcbqiZm2
OF+ntedTLxpGfNfUL+QU9Mz7TD2V3UAis5QBCASfIMaNG0MGCKZU9mbFnTpgAH4oh/y9wqWlsl2Z
7SYBlMGRW2pQ1pv++b1Fhy2LCtJ7UCvDdbFEIBP7KmqNEwSQXWy6cxAnELj24cY1GWfnOUqtBGIv
sOmZiA8oQz4GKS0uk8PJvIY9yPrEzG38NVEzmKZjuZnBKmjkdGDjylEzLfL8aK6g4fi+x0cCfizP
j15EWl7z/Zj1CfWfbJuh90WUnt9fCygSQ1BwKdtKd3W+7o01PUv+TEXqbSGyhhiRqLpjgm14mV4p
hoOswoxSNO0sQBkv+LDGurgto9So4xA2DSgALYugWC0Rx1lUsGFyFggtaaaE91VdIBk88zrI4Dja
1YxP82MgoXTg+y3hVDNRGl1aVZl0AEp9sAeh/QLdOTqW6Ge7j+jsvJBRnkdx/OI9nJpwaCWiS5ix
KmVPwhL8CY/6UDCGjK+TPvSrUkxGF78Hi4bQnnUUx9wLltrmO4YFamVJjB9EVDsBZbtMD4K0kseG
edUHRJ6hk6RhXBrtsNAKLd/EKDFmEkF3DXvtg91M15qXnJdR8eyMeBF4FVVHahlOBOGYgH5WwdL1
zJixoncQj3Ua0C4EE55cHwuTpNecSMCAaAA8bBarviSAZWGsgEdNc3PvfLa3oTwku1tB6idytx6O
Z2NdIYrB9ZJfoj+IePqee345MuucO9dRrjICFA64UkSggFybgsqJx23bvJMAGUu2JeDc7YCRGJIu
/cT+XxBEWjMj8HAjgqU8VRWjRgeElXlyRqbefVFSn4OkaDBE1r+ej2URlAjHYHLyykThqCDw86Ll
ipBAOV8eDxatHx09/QSsnY4n3aLG2Y4+EUYFRXj3f7YU5M1iJwcbbfr3ONBVF3EZGBqcp/iWjrSP
35w6bMSSLFmw9mPDuX5M6mfcjieohWssYveNSYHAu2fpwQAMB/YB8YJA3hl7RTuAauSOD+LyEj3D
sxCTyNOWx9DGv8UptU1QItji1qLL5LcWWUGSwc81bOlvRiu8KCq1fpOcl77cRyvQCodn/sdSipo8
XG+J7N193lnnjyvmIvYA+2QFtizrlfkY85QBxKlLlWEwczJHID3BOdrX+HL1bUKoACEeRFoBNSm+
XQjJfxGOtzucZ1jviSQhMOHCvGEJpuuMI90Wzids+6RI+mpw4kIjf0XOv2Qr8USUSHfzyKKw86fC
WD1P8TZXxH6uEpnQBc1d4rCYIGMoqE8uCwUdlvqUJ+Bmkc/tc3m3EzNc6iU54T46OvJKbjG9yY4H
GZYX1g8gRS3J1BgolPbig4YEDrmmNmvFP2Ec+h8pdqfzCEj+USO1VGB8xwuCeT+ua+C6KnhwEe7w
vMuVaUmLAtwUEfSHQw6yTGsDomwmVwYHhLaWFV4idVUS/xb7zFLQebMYBFR6TFbF8WqMaj2e9KXU
AV9ia8ZtPHQVS1ki7dI9tbPqHcYLso7hY1TipCcsGC3g3KQ3hXOvnbQMmGrn3FLOGdRjh5rxpOqP
YHxzhQYrlC1HfmsL41uXKaUMxsB17nWzmCxYofcIJGLBfhUf4pQEOf3Hm/rTEC+JLoJV6u0L4BkD
hbzxMQmrbjh3bb0X6PvzYmBekdH4IGm3UY+DzUg6hD4rdOL/bINfPXB9+7OpbQsXyXX7xh+BANFy
D+4vWxyN38ktOH+0DpZ096/qnyF6PrAw1eZ4GZRGKLmHBizCIdCSQbt4aPicZxYpF29ixlxD48Zz
tjGQciKSGVXCmWx7wUU8gJrWqSaD5mc6rXeWXDv+aHYzbUtlVvxEDRKtkyjD6k0A7mErFOLC5JER
+TiJvrZ2/eTGB7sf1M+UJOxCI182UN+RlfA8YpOm4/Gcy76ueUYrxfHacgmYlxwy5bIWQwE/J3lx
jeDhsm1sLofp3SOyZEFlVf06YFHZ9ReoZENXFQkyW+aQgntRGf7bLI/tkrx9Exu2ERNmhcZYnBeQ
Ettwm2RnnGtqU0r0A19/sFbBKQCdm3J/HgrPzJtvB+JYUoqnbuA4c1r3sYA7sFEFwKh40Qm5k3ki
DT/wtRSaZ22Jo4zp/nHL8m3vyoSWInx4H0aRGWyqxzjxbPccsEM+rmTImQbB653NS6fF7zRTj4FX
8MmdSBBqO6isdE0NbKJuvC19v8u2vCzhTrhjJbztGlozOx6oAVN7+u1VYVKgFTNnCewwEX5Y26mj
fdb0p4CPV7RY8C7pO7iNX98PvRVd8HWYlZ9uw3/Qz4/MnOfMtD32LLW5R/zqS3BNrwolhUvESed1
VgWAVe19DsJ5LeLqBhFcro665EAXVG/8E6id5ct2Y5gHONddDv5NmAXBy2rE02fLpBKAHwfF07Cc
KAbJatV9L+qKno6eU2/L9ts9X4HSc6A9HtblBjYTYh85zimrzBL9XWDTPp6W86APbPO+tfeaVCFe
tR8MbCANg29FpBE4jdP+slTa1zKCXXR4xYB8N55E5Q4hwkiMEskvcw9rqbCEDJazwxW5upRfnwNT
XfxE8D3QfGck7mYY4CEwUF+E64oMOVwXM5g4iOpEb7FoLU9H4anLrKlJ3463/qygfpFwhlYyBbLb
VbnDU0EvfusNTUtrkqbHPvyDRPOGR4kmifQgVAO4IyiRg98fgG8POnZsyID1OMiO8jcS2TK0qs+k
RVAYqBToX5cloWoiq90ZCobrsu70hnRTAVUhIRNaknRARK9XSMoEPxybwA8f0spwCUXv1wU0SVrB
H6G5VwVIh9Hsa2Yg/iurUDAs4NJ8jdxlyOqu/nieyK0eDnMhOsjQNZ0AsRl84PVNmyZcZeuldETY
KAZWpej2x23Kmd9iPgrhtqsa8aykibGPUFFLMR4WcbatyVEC9DLxzzSEtfzUp4wct2824Knp18M5
lEnehoKaMwUNu9VZFMPtdG0rDYM1bv5OrKaBLyoQ/rqbgz7g5GDcsv1DY+e86C/2G9pQAkezOkCp
ei5u9snkvrNO2M9AbjQB1024v9SXblgQn58eXDupQeipifYd6e+j6X2dJHO4Yh0OpUQ0znrPe9ng
9+eGQDmRFY8EpR4bZ9362wKeX/U77BfVxu1lFrWKZze0M/VfDqUL/1xHFC7rGcJbxIDsI4ABZVdR
XyiQFjDX5AcKWKg2mZtOV23bA2JxYsby9ZXpLvVD0qcH1QV3YXKPcgpuVBpCqvIShCmZ43fgL6io
wXPRDhE0O5n7WBAilhW/aX4hcH4du0KEPA3r6IvFvLP0FyIW27cHt0/8WqkbIIeisQUyZP4KL8Ie
m0Tmrtba3I6a2qLUg93aHsoflCCfZt+mW1LHYf80wKzkDfNNzcVZraCITlTM3Sckm+4Q1vHemCRy
xhe920tZqdQYzqB7N+/kHTXeIvVVrE2xotWkJPpBS2CO8kX7cbFmY8MOgJ+OuDBtf10G4wDgC04V
vab08t+4GNwBSLPZ9LB+KtXGfBawsS4Rfmkgv3/TBSnsJEGKGLgcC+S6M7CkHmh4ZFfHsRaTilFW
X3+Uz4HuD7egHrHJDJpN08cShwLWpkdK4e6dH7J588bbUH8fHdjZ4T9QhF7QFed8bb39oqxBx1sV
KiZUOSd3X+OzAMo+vNbqTX68OhToOC8HzXhLFz97SqyrOH81lcm3Jyo+zn9BsqMNKn4RQV07jld3
gAfAYy43RQdLFM4OT0BZaPmblFBKaR+qyI6F7PhigCBk+RHlKJDCSI1pE6sWPOKE3P0yPjdRuSnX
ZMgbEWaRWdfPocRz+OzeaRHUHZB+vvmn939R1Ujo3r9ArQ6KM3hX+If4avF2ns21IVHA6+XAvmPp
UUz0my2I7elX8g1Dk+YEJRPISMQlz2CL6RGdd/1QmBeuk/1xPcHz5a8XTl5kiUYRg+kzXRIk5KVB
ItvTHPPY8nL3b9XSoBHmbihMdJm+I56dvmB8jpDhh0qvAva9qAjSJBYED3cYq4wDebenmW8rIbIQ
LLgvlE+TWZxz0YnudGsuVIs8zCYFC5DxNpwodWXc2v4BFI3Jmg3XBlSIAsBlVNw0PI8MTZcXRgTP
orZ8+bs8xktTiy6OlFzUJYhR14OWJZv6peDWlN7eVUrsgMe5mfo2/qRAzDvBNQ5x7T9WMJhFDiJc
HKOKfMElGDpmQNb63jY30bj4miIZxQvqG06sX7ay4YONhIYO7mO/pp3D1i2ccrpP2FI5TqHl960V
Aw1JVBthitx3KH4qwsyvoT2nNizyJBhfh9wo4mxa6wPEi8DWJcqmq5FeZM3AmFnhPn2+UgpgX/wz
XTCKwv1lNbPw8udphfnLZ0PiW4BWtyFRF+m2qsI9NvsitPa4OqApFPAdbDbewFzheDFGq8rv8Iwt
tjqxAv6VARcQeTyoNCvJ/Up5Bh/KxU+FUzXSNEKz7dGE45Gb6KvhaUp1xt8yl0gRVlF99P+LJDF8
T2ZK2TPKjLV6CZEtIav6ytpDMvkDB4nRyTqMDX26WAWP0f/bvuSvk/ULJ1lsAQjuFzsB4G2JBq35
P1JY1EoxwG+yJS875uYQqOXmffO6I656Tlei2S+XOIMMCSnpgf6S1J8mNw7jaJFs8ZTPNxmHU2A0
uM428OgNHnq4+Of7r9lJkfj0jz96OrTJVPDOGvLlSNtnQ7wIHujRkng5ih9XpMnURMsKaLo9qiH/
v8QcwMV/dpgu7O4Q/pva7V6Nx2qd+JlEB1JtKqS73J9mptMkRjNQUGKAvrIng7Cwn5PLEWip7653
BAApM96Z5c9V9fSt9uLi20K9q072ptdS+2SU4tbkOdJ0kayc8a2uS1zjeceGBfbkgZ0yAEFcfb2G
/1HNQXYBQCrB3KL9fBdjz4wHp/AOJiVxAFpKq+FlQJqoTuIqdVVeNzrrYzjcV0LEnMBr0IA2h8et
Uy663i9D2M3minSrZiZ5UtNAFkp+z2wUvhOIuMZ1fLA1SpxwqPmvUdauYoUd0m48FaJkTwAbDcY+
TZAXE7wH176/hNVEcdAS+yBaIwRTpuSxX2C3/H48zfOSIBqeE5QGk3QZY264V6gX8gH7mQPUaFK+
6cb3cteP6evb0CPcNxgaWsym7BZmgDzl61V9GRAaXt2p5bADF5G0MKOzrVS8AonZkdjk3WA9uFjC
ZFl4DIadT8WTA6fPdLOnmX7iIb3ctaNCtAaQgqF0V7qec+lc6gqy/RCdV9zQ+FOsOZG7LMjt6MS2
8tGYcFibYQe+DEpDZV4cR+DT4Xa/Zw4Q7uEPTaypmFL2dPQNyfWS+W6JTipalEc3ggf5HwDZMdfS
mjgLcm9CdDJ4WA9hB0edKsktouQO3lb5tnchIwXNlR0T0lBjIKMLlXWI7N1vnkSo/ZF+WcF1iNPo
tIlexrMDLwan479lVCk6rL/jOXPQ8Je2ukeOCFjvzegQNYEIt7GdWtYZWPQ1bk/vkgIDYW2+4omY
me6ce6tNizuc05rNwgZmEylLgIc3z41hrbGVHAfzRPZMJoTv+YBYc7hQUR4U5/cdtkrXRlY3C9/e
87sDRfPsCprJXXJooQLIoSgdxQCTQZ4rIHmeyEtc+FqMUSR8lFrMTXw8wYUsmtlOAV97bO+DpJr/
RAvs7uwAereR13G5HCxIFGzmVZ7WaJ3TCP3Ite1BWa3wsO4T4k/9lq1obzVYrFmFgv59qDmcNVU4
YhblymOcd51EFFYdalmbWenzboF4FPZF+ULj2gmLBB+980X9MR4Yok6M5zb7j1PfZahI5wtSS5qB
yHm12EgkbpTTlLIC//+Tthcr3k3mE58bLqRCxGzk6J3eMAug9Mwd90ZnPbi5/zEiBD8WXWhxXY9L
laCUvK6vaQgjYnbXAkQN7xkXynuxkWR+zmlwa+5NaVEvFbnOFAJ2j+HpkBmtjYTMdLc8MN44Bswk
qE/gJEhqXI7XpYcW484LtJN29cZ8SpRND36SFPNZsVUWul4kLEHrAppKoky7A+FtCjjr7srbCtmC
m94cymfjWeVjvyG94hDA10MVElvg+cLLOvqVsjUqRKOXIqrhlBEzehtG+NbyXLijrz+D4xtTw7OU
OOlQo1wVtmhrw9tXow941Wtl2JjjUFfkwE/KKbjg8I44aEZT8nJNYCpzTS1Ceg5+z0j2DN92KzK2
hu5Z1g1JvHTx282O60gorwyJPIZAtdeUYOujhMzkS2aUDOzUicggT/leyYy8NzKlLzHn9j/nCXEI
oZWOoCvxER9IkM41ebfW87p1H/Y1AXGI5Ize17S+aue6JdoDK2nQsbVDjIE+mgDHCsW45ENNd8B3
U4D8iHA8mo5g2jx+DmVw57ArBmNGWKxhIEKOIAzNvKW54mwn1rylIfYQLaNnSMuaDlFUUI7i2NH4
9AIvObN5ffo+GRNFqYmziJFc0ihxCUhJNiAlxd4M91ejnRGMkOX7iAlULiXdHUA5F6Y3JFLYRXpB
dUhGhHz0idl8OW5yjUWYOSkMgSUcjH0cd912BHa41Z9gmWNuYt5CwOVFDTKZ1QClx3+jcpBYx4mS
uJdYqYjzfs2ybgRPn2C1EzL1KUC1qo0rGeGQFzDEPBY4dxU2GsA2kFBZaiUOXcuTt6KuWBsKpCbn
8sq6tAlw1EMg8LN9J1R4fG4xl/cIXlnYkIVKkS6DJITpp7Z89bkjMngtM626zLpFgoUUocf3UoTH
QT7GxNn62PtrcX7rbrMbuTMtdmI40IAwVbVaVHi+N5Vvk8oocnDcBxBOdCMLmc2uquMQv56Liias
i8RoWFNEQfyO/TdVBAo7UFKItC0y46JTH9jj/KOSXpt00PNx4spKHEJsZv5I2RvCPrQ3xIkofMvD
jLs4erflOSAk3jqdG2o7D1mFrCeY9ROGxO6y0whO6e6KvuO5hUkFb8REzbmOkKGSooTC9F4Y2Szg
qixgsr3DSPrOXc+gZEinsc1b4ZJM9W+WKA8aW/RModtU3bNSrLkdG1LMUvb4nShJ/4Nyf1m53aW0
RiCzXnepTibPId6/uUJ+VRekb2gnSSVW1k4X02s/Bn2F0LRp3ekZTfQXWM4+eIocTPwclFSdrzXK
5YKx63/vytXaPitrXeLDCYQ6m5PTi5A5UaKlUMMZ1lfwlUBW2dcCXRXmNVqu8pTbjmgF31/i18Nx
sExGgRPsq0CD9GBuJSiSGHhnY4Re7UtCqUUY9xD4GQbxmiMOwEvF5Xo7pQUWjTAxmaXwTEciQqY/
JW0Vc+FnqRHyLxCsx2XH1orRWozVqRVw4MmCm9rRue9db81aQq0i2a+8LnMUi8C/YOKZ7NJFKbol
qwKnF14utSow8gzvZNSACkzcv6TacPcccm/U1yJtn+vdrSbuMvtkpX3bMaaaMqwXpMZ++1oFG40d
Yh7VH5GtNlRckMLpChwVrQjYwIQNOrSD43zfpHMyWXfAtcQKDJOp1zToeSO768semwMPRElmQtsB
SarUyrXHL3RiIvZzpotwFKfrV7ifWBy6GBLvW7fTulG840/d8zj9cSZO5q029JHDqbCiXlAaY/aQ
w/zGeey42CVJ9iZWWfzxzFbzL5K6j3zyGCGET5Kb4s+L/uSDrrln2Eb1B5Fw2czBE6vrxXTdbVXv
kny8LZm0v7RwhBFQvPYMzWfaIcRYW5IoqstroivCq8Fo6RbXEXIBD/a+UNgNPRJtwx7o3ZpXfgPd
tFfxBeCXd1FH/0KCGFOsaEsm2ZjlpoqWfqhx6N9SoC6qRl5qABheapi4Uo34vUPJ8BUEBxiD5UO6
8upsrxiYfrdQ1h2FvvZEq2EkZvah5QuRzsoV5SoA8KYmHs9DKj1Dog+M/Qr9qFMGGOFZY0DXes0B
AdCUIBJ3yBh3mDMPdSPSuZvoKDuynsfx4XaTAjiN97f1Muu8HifCJQAFgGt30dowPYenRXthBSW+
GuUvNyQXI0olSG53ohlMRpjy89q0kOjEuI0hvZh19yZc+gdDiyNvZ4Vbi9R9DjstPquudigvQiqC
S07lNgbM1v5QdVUc+Pdm/MEePSul64+5jYQRF3hWnR2zVLFynLLo8CQVC4QFlB38OuKyN8usgHSn
tIxFucEikb9bU6ZFkwhuiffS5YTvvyRRbEWSTOkGdsgTHEmCMEO4mRoywu0RuMM76hbTqurHDBLp
Qp3xAM+F1cJ9dToZ4pjXvnxjsuHtotbFQYgdzDW95imFRomE84VDFvobrC7ErYuqRHh612R8kglf
jhF0oXLjpF+j9NVpsARk+Gx+lowWpkj7s54M2X4GhMOh/a/VIomzjmk+9EnvCgEAn44LjusSauR/
zPv/JIbRJPTX3dKG08n2hH5gsqt3LcO8K36jvAcNDgDf8aIUFkkLx8iXC7BQ0riL5NT5WRLqvjr2
TKusemgdlsbvVLAczyTxNtpwNmcNJcgCJbXHGMuolxL8V5npPgotMqKpwJFUeE6mUhi6U/GeSmZw
8mRu4QKoh63DtS0JmMyYkl9Ej3jRo3fDmEyVU2LO1TbYO2RCXxQMSDPHXMzIlwyd2I/7s7h7ZgM/
2h91ekrj+44E35rAvyVWqeuskKQTWyrTvv021a1cZsZfoGYyX2BqpWu8b6ZKDP0Ry7Pyu02n/cbE
s2W+Nrs5eU14wz6r3Nkmvp7cxbYGsAub3CjW0f8K+hfoIjArAf9NzI4kzSGelGr/MOdsJYWBy72o
RaO2xyLKmpHPaMQYJ26PSl5VW3KYWUGi4jl9iTDYlcu96e53HkJUPPMCrW5HMoSw/vfdo6Pwb0gv
RqoA9bqTgm+w1ShwgdXR3H+aVZnghDV8gzkDCRusarXz2Gc0blqIolWOkP1veoAcF4Vuq1GOTCun
gh1w85Ummj2QKCCkGU1nv/GmtVSEwOkiuBAeNi/MBfpYA0zAKLQnFbhmEjNH+bBDPOq1MD54iA3W
Rvvr+gCIF4tuA5R9oLJ9ux8NcZzK2R4scqshI1HskQdMiNq4FUFI702ncnGf8lr/IMzMxs/LBo+F
Rt6Zp0v8x1xHSU75Dy4m8XPJ53nowgPJEFW9ZX00M1GYmwczuz4uf4oQ1dR0KxwMB7LsVuu0HvIm
ETZs4Pq4F/Gkdw5GBzkFN2WjQq1LbGWyDSkZFfm/GSSCwQFmx0UqDkATUhLVMt0emivLi2sz6WYu
WAhvuY9OIXSGVFgoxuQ8ZrCFOjQ0QhrSBPh7IAolJPMUvkXiMoAVRIjGz6NhqEFgHX1fU1Drt2UA
i3lqkHLLdRTGffd0hIBHtDD4ajQ81Nc8ADyEyoZAKSL8D9YZ9gXxdXzucwJU5C9u7eVKbb+a3tmN
PC/cb5ZutneYeM9ckO+ZXtK+Yr1bb+Taddxj2vYXcaQPblqBH7YTgYeXcV7f3QEb45RE7noQav4F
8DHY2dI8fjt7pq2TGrpCNH+AO16rxh/v1KPcSd6P97AwyNjrGYSva5M1iEpNwbKQC8QzKIxcVFSm
Nfw1EghTMOjAJh+aFF/7+DaHiur2EpYLvN4EEMgEdDsUoLAICONsqErUdJfCFPFj+DxiG1gDxOqO
/S4BEt5Yvm+h+gl3/Xlx6dXC3VQq/gBcRG5RcOGHEG/YZqIpsCeC2gZZmD99Uhfa2jJg40wSWKQj
alMtZH6joKY8ME59ycVP/7YilDYzfprye1Yh9yIBnJxsjaJrQRbXA4F6vyoxLgYaHpntAuLw8wbn
HugDG5LUq3dmSdYryohLCLXIPDpZCF1Z4UT8No4lKRaHmqw4yj56e4DS14K0U997o+It52YJo/EQ
vieWMl9oFCpNSjm+YmZ3MGkiZklDTRxhWDkU8VkYWKVLDR4PBXzsKpveVlQREwG7aiMvzN++qdDF
ikGOsajQnjdEh+poaeVaqAeEeUErwCaXoijG3ih1JimHU4IgHcjSj6dQht51pPrazVwl+bcGv+rn
UQIFDLumTs2gJHaeF/tq+G36/PFiiXhUEE89dIcxdgDCtOkpx3RvmihtU2tyDzHRavj6pJlYrW6C
JVJbJRS0LbhEMgjvzQ4mgH7dGYgO1c8m166HdeWST0gFSTEDEKCweukTzbtNT9r9DbjwDov5qApw
9hSFDFCGXANnMDxbEK7HVv5weDAy1MH22OXxDE3o4vm64QaRB6R3yQMNXFHQwjLjz98Gzf7JSIFQ
mhHrkM5bq8kJp7UarJemP/hS1b7XqNrUyBrnRvN/ViE85D4CIDkaxivgnzFucpS8AijU1uL7pZ24
5d0gV+LJvBwwqjoTw7J5FS+6o8dlg3LQ5oeaJP5RT/izo9VBMcqSs9JtI7t9IO5PWv2M4lb1rJie
SFI4vVJngsFLf1bwT/rFbO2ryY3XZhv4gzUxKkzmv7x4P7mF9WdiQVDrFEHqahK7XE11puUZ63TU
99i/4eiBY2+cHMIBIAUZL4z/oYNgYXtNEeSjACmjVJ2+/EFfCre9b4Q1Ih5uD0EicGqjEHgjOzFz
fFoV2QFYdxg1+EHQm/nf+JZf1GU9OLhvuqo23xEW5ctdP7G5xtg6Fi/+n8dpRcfc/cAVDdOxD5nR
HTYIDB591jlvqGREn9nVdSVxFS9eYSw1P1v5kilaHV2tgP0smqD7PNv6iavSdAu/iCJPcjMtDL2x
92AeS1Rd9B+5W0nWZcs0mZYWp9sTlJ0Tb9oGG3GmhMsXcskUEm49FoVds5YKlSm4oHdGXN/hP42W
IIjF3DBnv+YgzdY3q4UZTnt1m0j0szMlvKMV5hMU5UXKme486gerjD7N/1JxfD+t1JoBX1eNZNwq
80pnHQkHWwG42wSEbays6Q1MS3Al+ql+EM0eSr3h2niKF1n9e3REfp7VOb0dC4wetv2felTh5SqQ
l5aNGm3ExNxuw41/jB0aK4pR9Jy91VrRpyf60eWfjLWUa6gcc2oien7UnapFhTlazW47VKhAl1dk
xc+sdbSH7/eTd2oS4dXEFCtFIBbWxFnnVSJciG/QoArAcR/RJ6KB0EN3JY3ILZrlOr0E3KXZ9EWH
ZzNvm8dkXvU0GR4lyTRH2Uy8tvzP7/ZBsnP8x2hGKb/gJWWPSq90kmVOyWu5dArS8/GFEXJMOevP
z8UJBZ1V2Ck03nNVG/iBYcsbCLNyHLT5o776Xpfss1/+yotKbjbI5loGcNRdVtkLouratZD0QmkT
bYw+V8Ro43j69caWnIJZHkABZPvf9YbhaoMuiS5CAlZBUTfHokKtvUj0Fe4eeC9N1n0dRjB1/S+z
OY3sOJ43dXVbywNd+W7pjnoay4K2JnxfYT5yTqmEzyvazKV7Oa45a80Afi0k7zdiUIteS+RQnQT2
ALkXT0l0562Dnf0uwSxePJfU9OCDhd0lrMjqH+7XhLOkFzXrvAVPx587XJhO/ARFV6ihMLgedq/N
R7n6Xme99l1k7Hhta34FMlI+Qd7tA1t35E0m542HUW9fdRuExZCeKAkGdzT4vvw8J5u9wZKs3IyB
L/o/HWxL/k5lF/nAv6lY35uVwUH66NaLmSh2aRhfzJn4GCZnJrp+Nf0u9+wKBnJJw1FqU/wHhn8Q
91015T4X59ix7b0qL6HoOCPd9sX6mxcLLVUfRn+54qNtxHw4JrDpj/Ok2X1pGqfaUdtG6JvoG6z6
nx5xZwW98oUX3uIzS0vV0kBVRTL01NgryXdN4qD3JIUfCOwPOtYy03aFarV9VZ/ReQKBdLB6RBhS
zgzQNFyrcx+5HPaRGITlncyH+Ejy2PMokaYFf6nLAHQzUHcIlQXk8w0beI5K0EX9b2qP3usMzxrU
88wTKfw2R1EiH7NIf7F+fG0zf4f0Iqq3U7kMU7joZNJL3UwZQXjcwXRBqtm0QeCZ/UOidWj0exFL
g2KI/ar7w50Hng4R38YFlnpsDT8Ig2SAZccg+pvgeX65Sw8gR7XLetlwBV1nWokXAs47aC/jJ9h+
i+QlF/x0RN+9BefmjxtwzJN7NrqCzFYuW384qwbxiShHEujEDcYENy4ZeALSUxPOAyfm9JQt/sZX
N+BAO5AEXJ4yGgZtAk22He81IYjaU2sopunGlXuLwNcs8C/5Z216OuebGLIaKMzTNF6SX0jGySFC
O+t3fC3wlqRrMPWvMqU3HHG2+EahR9BDqaqLSBwCSSi0mkCUUwS6nJ9B9INHqWGd0HXg2ERpd61q
gfrSocsoX3FLz0Hs6/acIR2M9nsapDuJnORbnN4RduEgMXc3ZiFrByw14wx7SjLHNcHT3L3Y+qFs
luXmRnp39CNxkI08pSiw6oUUtybqpT002rwYnIDhxaIhDdv6aF6/JQ8HNXju2Aj01FxO5APRPMch
6kc25Tyf5rzXNZTdGRV2AVPVWUpGVRB3Z3mD+L2OZ8SH+kSIDdmH0Mo457dqr2SiHYcNoKMCNVVL
hqF9eJ9KNUNf6f1fpfEUFaSWQ6h1Ezllw5R0LF2+TbrFaxCa3Bv4C2xmk34UP+d3rtQv4O/XICWE
Q8ddeR41BHx0pS3ZOh0xVYljdnZA8cd0JGL8oNiLPWu4PD38x2E0Tzh/h4th3uVZg6107kXQ1A33
739hBnkmRSbxjx8g7RpulzaxJ5CXDFiKNFc/27fxOR5T6/P/4bueb0MTcyVzxUO56XIXNF6XeuCF
vuKLLhkrOK7W2Kj/z09/7RkdBhQCL7Ev3qnIKjkc1nAE4Py6C0w84xySVtYfUxum49Y+TsrtY2po
L16UtJS8ix+Xn9MRxqn84YddlEj2ht00rZCHWt6DSEoUhLBYORwApONiN3ILHxEZcQJqyJx5cbNk
9lIkxwFmQnQ1xJ65HbnWy17EDor0FfvWDzyQqZy4jdIWuTLFloX8hixP5w4ionxR+Ijo6V0/3W7n
t7oPlIGneJBXUWCZS6KwqinJ+kDnlErHo/1Kaagoi5wMXUQysfE9N+/G0iLmCtqKsWd901FSxUuf
OXUROF8NWE7Z4Ef0LScw/7d3SgXeE85rys13NCeIE8CYHIx3fB6KCy5+w+lqQ9kLEf62FgIqJB/S
ZmwJqVApsNW75hlBjlyhVo52TtNq2a1gbf0QupypOv66OFE8KLtoFnxGiBfVruIqGQz5LisSfBkd
7Jx3MPJT6Y7M1voYXAWAK/8RPmh6K1quM3biHK/gFbScATrsdtueDe6subJC4pThtUrx/yC5dTBl
LbpuccJetced2v11SyuVp7FAbyPsv3t+w3ysvZrJGWUgw4/bmlvnbecX+I3Jf+psgXR8nXdqAuai
CkStGK8oqEv6c3IBG8urqd1lbx8wqJvxgtMoBYx9vNIaysLYC1K4tUaFpEpqotwd6/lXL0Trm3bo
1jDxUikZQYOEvyWlmkTJShceypIbUZeRLZahc7ODvCmcvCYDncbeoMoK7Kwch8R5n5vhFoRThcOo
3SflgcJQ+25usho9siLJ42Uy0uy+dGPcnOHoUZBASXq/TZhgSZdjDShHGN5FTI0OtEQ3QZDtjv9p
ymgYlKFmHfwEb61MVF8pI5+TW4UgXNbt50mAKIPk4G8dlupEC5BYIb2CRW5Jo0UigSpJ0rvw4MuA
U3pTK90BgyGBd6ICdseMJhJopaXXPrk5z1vu2KnHcKvqFKNgJ9PRTRpe2Ln4h5E/Tw9NLeuOzGNX
v2g59lFIhSksxEo8z1ebWD1madCBFQEMW+SeZsssyJDEqzmCnGh/ntos3A4vqAW11WGdvXCzqBIs
sWf3yJFC4i7mJbSePV0e3bvGQu4ybjz6VNYFQ+ttyez4WryeNR6nmy4Vw70iGC6LlInSds5Qs+pa
Thcky48jU7OSKWynio53hTC6IBgcG4jIqnIHAsYotIBJuTtXtp8RoEv/Zj2azF5Zbvr4G/0xF09Y
+EfkeffzwpF5PzQrR9HP5SM01OenL6GQiut6xJTrOcG3BI5dLBkT7a67diRuxM7qoOOSAcygjU72
8bpKzBhi2cXbvRWfTmsqtfU0pxn2AZt+4EbI2qxGQuTo/849Ih7nc+yiYbPxmqDnwL8NTVbHgdm4
nRklVR1jpTxgsB4p8DyOOYVMcbwDuK7YnGFXGDA5bkpzpvGZWC9d2Y0oz5fPRPLBdd1124924kfy
NnS/J7rSDIAi0ZuYBptkunCNl/q2fsQix0uIMJF9XUg0+y7SAnA6W/pVMglzprxkf85nad6zhdBS
SwAuLhK1Qtvo+LJXPhroiIvbtjCXlCsYSu6J8aN9RdonZzK/fs3cgEYtBfjIiRiWrcf1N7lKbZ/K
+m2PjTfEky4a2toiMlmOs/VsyWxzgEbzqZ+ARZyzzdmvkL2WqHkzcntGHHNxkMJf4uu8bOJbOdtM
pqRJ1g/Q2LY7GCwBMmZLvRfFfwaqR4CcuxQaGdjWVfl1XykKxzv4bFJOnB921e9Qqi9il6B6zuZD
3gVuXsEENA4YxEwYTYdMknfZ+09gARdB/YE7k2eWW4QpDEhMIiC0rJmpok4YxADBfLCLdBffkN2j
iAZ13Kn7o0zr3DvGTYzyRvrkg0LhQDz1o0jc9PLyuh9QTpdtb8KFXwaUmdd+bND3OrjJUGcHAoYC
f6aoHoC3KHVVYRocs76rVGA0XOIjhDXbhjdcouQYwkXGCQcBjS5M4MjtirsJ5m2dP0keR3tUHX80
sve5yhePZ25W32gIeUuE0EEpINiiFK/qGYWnGdv3xMOiTEg/wgvMgCzn/jt1yU7f1RTJqfTRO4yH
APr05XN8/nLF6DsWBAbyjaRseJ4MjNZI+ulmIDXw00JCR+b3boSRnxqMc5Q2GgS3ufEMzBB6f40p
JstcQ3/ccouExe0OK2Yg6TwMfU2jA2fre20lkYQRIceAJ5JDI5aBsBWShx7ZTWzpsSISY/lkJ7NA
30QEbdK0pevbQbTnpA+L1zitaSXp1P8ow0a2IjWfe6Bt2TSXzQvRAqYFfb6XFaqHAJihzSMB7Ub7
m/nHmBclnIs57zDAz2l9nPg0CdBAt1y57UpDDPTSpZ64cdLd2ITPgi4TesptIuizgX7fBWNqBJp2
fn+QSc2OX1Xa2CmGn+68UVZL97qbMryROEb9prjVu+sx1HbkD7MhumJnHWyHwjR9VMRnHHiRewTD
kJuEqfcBm7cm7MAcGr5/laditdoXIZZ6lYjmnHxch/uPmKfUdA54bTCzFjfS0wG37PWbq8oa1M08
PZNidZrwRTXP7niKEJbVfP1dLJsvLcdaQsjMs8maqpWBbMoQyv4HbGnHT+Js2/rW2w4Cke81E0rG
/79+HT0oHZlqhgjSimsam4qcAZhkpalTR/hTt9LxlCKEzCCpTVRkR3d3YgKnSrOW6aUPDUVr7RZ8
rPY2HrCF33ZmSAuRPnGGWnhwMB9YnuvrGxKh+NNh7pWOYIwjMr/useBZoyqUmC4jrdj0ba1Ifu3L
qhau4ivnZ9fdck5KfctmjJCX4snVT/arcwIF73oP2e6MccUap5NQtoTXEaBp8ZoqFsAuuyPTSElX
ZUKFmIjh4fjO2D0TgBleuKOqYGo4tBgN0AuMTOUzYszHqmeId6EBJJ32FjT3drKN+BmURmmDQZb0
TA0hy6CtKgBx8CUG6r7bwFR0YQZMVxucmj62IJ0aVOVEhzF9aJuSwXdQKx1jOVVzOniKyKjJTTqA
zCphoMzxAk8BiO5ldrgU6T2gHRcOt9x0tFuJG2J4FHdQlf6mcZosivEOGsnM0qZL45PK8AFlnf92
OGrBjFEzSGIkVNu82wUnA03Bm1QqrbtvXpMej1/R08PPXbz7QZh7ug9tR7986L+jS190yuM20N+T
2CukXRW0tE1ExrirDMBqu5Rk+C2UhA8f8ExQiX5IQedOFXFpVb/k8r7KipMah4A81hcRvEekv/Bi
5Cck4O1V7a+lkeyjUF0/mMkWGpvNvn7XPe3gjfqINv3feZiigbt/M+cK9p93A2B7kGpVN982Din0
2vIzW7EyhDXKCHxxfg0K2YiATo5hyry7AjSXfAtfRwLjUbl+a9PtOHbiOJIDcC0XL0Tsxrh3X/sG
KROrxZiofs8DGOd50dokEqzahi/kpctIh93A7moDn2AU95uzSBNUNx9+K2UAV5eI4cMdPqlPdW9f
WYcr6LyUqmaApsadtLv7dV5zKChfumF1sj12SHcfb1wy/0jAd5EJ/gjRndf7nE7l5HWZ9ZyycAb3
grMn5G9sqK0rJ+/dySF1nVOzoniPTeRGxeZ2OTjFaoV2qIllQKuG2Pp10I4EGvjQubzVgHJflpm/
lmFHxZ2+7E/gpon2BhkjMtQ64P4gtLS1waUpiqcFK8j2NrJr6yuoEnkPsbFZDmp4USiKQtp3B2je
9laCTw9owPP4X2YuQalNE38PmCCDdGSIBH1wIWjnHB0YO26saLcZ0cmJpDpD1WA4SJbEIOCndsrg
MtCfyBBXfyUsh4srbggsOb/0CU/48+xNgsTGmSlwqrWC7qPh4tvxgZB7w0LTX5mtBrMz8sKV5BXx
giCIulGa7kJ71Stzblh1bgmTED16v5rLklNrX2R+FCyimSIBiYLKgaTSVTOLwmRn42UObge0+a9/
AjN1jw3nSysgHBkx6LYz8g6wB1jnSiT+A0pTwXJDUiKnbniXd50DI4Vf283K5EuR1oFE4P796ly8
iINBpNhT0AAdOJoQ+X8VGXtv1B6VDAaq4nYiaby/AC0BF3HaHGOblBcl56wDjhwop5IemzqPUgDQ
biLokBHle1vur+fhRVHBy+iwnY43xyV0HLo631pmAbiZ7581yh3E3NRE8/pQER1z3I0ikK13x5d4
A88a9V8JfalpM/4lrsy1RxMzkrG5yp7cWQAEi+yI/pokQD1bL+wG1BwxprTMAMypGY6YTwJ0JNVC
DM30+IC0BGrVIz4j27BnF/zzPgWXubFMW7c8DwermUkZVPHnsseDeNGI56O262EYBAhE4cuxLTVh
D7vcx6+QBC7AVRmiYvWPRlkrbBPtti1u08X9gnhCrUXYZ+6fizE85LK/BuR4r4tnCvWBEG5VuJV8
Y/j2sbFaO8Y1HU29V6z4Nl5/maBgOc2/+PHdTNcstpO7ccQGHJrBonoBaaWK+4yf/LBL0wp9FMNz
C2xKgbk3+4QODAeiIUcKtk3sgnQ7U0vuMdqfNsJEE5v8FbZ7IyZx0+UURAIEB2e3chOF9jL/xJ2i
VYulG4JteM2M3vak+FoI8MxIQuu2K6GDvsv1YZm7OhXyBZsVU8+8dw6x2tJaCTerO6KjTC2zcGFP
d3rUSZVWtv7TYOn3MmYdhKmfj5GuljN8Sqq76viXIlzlMFM8/ubcgTxW0UD8b7tPuktwSfG62s+5
vTek6q0ui0FnXfTHHnrn1KD87qY1GGDC0S2iFVvPUkt89cgy6bbylS1ujY6HlzouewcgkrSCqSDT
5TKtP7A/JQZw/OpMRLpY+ebKnP5LMVjPeCsmdED9G4TH0yhsrNtzTFPErZxvQOcazTEnlkTaY2Xl
yDGiuWx2unNApEJG+eVNt1yWxmzd7kVDPoCFHIOnZyrUrEwk5mROtJ2tesd5M/nPAReelkvMBgrO
IAmnzGh6UdYY4QyrrhxXFqWhQJUFoHP6vM8YqGbhAqz08yyVvNSHjMgUeSOmvezikjz6HIOIxABW
Mw4wMQAD3dJDVT/WAc6xzSwvHTT/cleg6D8n+MG6XEftwZcXJQwyKC2LqxgqvNMfwED7uGhuGUTy
jhPHWPVB+W2EWWU/mWu3751HZp5Evb+HcwP8SIcZSaE/5MwDn25vTSjyfpVk8r8ntPMjvtQWK9A9
S0AUzBQRJmgawK0usGdUyZX8pJxs0KU0XM3PEPMM6qdmR5s8hIFU83hPPv9tGNsEm7e8C5U90dpe
efX0Ee1PWe1IfVder5845ezlWXKl1WhL+niD4LoDqwoA071uJ8Wys5fOmUBxrVISKFJlpZaesxxk
qgc239c7w7MAn5jrs+4JHS8WN7VasyKswD0E0IQb7vd/k4bhdO3TEm3BQkJJnOpikEuhUA6FYVNv
1V3wJdcyjHi5Wo7KdY0b5uBWjCrhgSOQvgikeXpndDInnsznNkHgCKpxs9kfIaDIv89od4+7c/mb
9MRuWr6vC/mdbjTFZKYHPMtM+FE1vX81DtEnc555c2UO7X6SCR8Cwj6QBY0VfBYvaeWDHChgnSyU
FHBKIsQvSFPZvK1j6j4BlDnAFeWT66n7CSmuh972TJkrw2TV//v5m/AL5m5hkbRn1HOwWuVwjhjf
VDfeI5DO01t3WqZf/0FXwL2ciSw1CF5fgjl8oTHB4BpfMI1Gs0tB8d1lJNMQSi4iWoPCbzo8VM6v
TW73QSrvufRZs4Zk6VEdnwAUyf4uX5IR/gfCTecwMbn6NA2tbEGkBWzu+mI6h2am7/MkgPQ/uTVi
VfJuvIkqFq7DsxFsn0nxmPGfsq4FH1IFt+f/jNCTe9ngR6wmt5ubaAtAFuSZKujSvT+s0JYdb5bP
YIJnj4g8PXHoXD+1qO+4LzsbbLoaD0ncJalW3TMEcEzsSlq0B5pge4Y0qAphsix/0yNe3wShESvr
fu+tPSd0Gwfcu0mG0PTST1Vv44tTXPJG+SRieXaQMb2+/oDFoYlgkt0vhTV+xeM280E5tcd+VkCK
7jC3qE1aO2ChQT3NSzYce3aSS3JfT8nswYXzpzJXHvk6xBekVeUBkx6ljF+FvJXTFQJXj9hKfVgl
JimUIbNRukj+IOJhKMuOXANrR88fN5CXXDlF8TkjcLa8VctjlUs1fWyy0yJK6rwND0KthoL916Pu
vJBgXsoDq5Cs5oad9aqCJHyHLYe/fen/RBwO5yFrKOVqTnIz8gb6/h2Bctfjl/xM5DAUZyJrRtlD
pnjcdzzQ97ZlySSiyof31mVgJYgMo5vnAs+UotwnLzO4JzNLcvc4DF5wVsjk+nQz0aeDYKqX6LUZ
OWnKLzNqhXF9YJJ9waaBcTAanWZrihv0uvnTM7GLwtjONvStj/qy7Vg1H9zIP2w0tzbdNIwzzgR7
IxQqi6xYpicWa5RlrX3dRhZoWE/XgS5Zu8aQOiiMF9Id8sNr9jyC1OjTes25mp5yoeiew71x2ZSg
2GIgDnQ64zZbIF63p7imDV9GhycdqcdMOwgIjU9C5ephSdnhrnT53ZHX0gjJNkDlJRI3vrNYCsr1
d+TjkGbgRBOMs8pdYQP6xsGJZvl92X+5Ec4yi3kzinc2LFXn8tGqxX7bqSHNWxptzfjDjUos7G0+
KBQfoci1/KaRttIvMRnGKUqAwtu9ZlNIYLMGesq2EmK7xWrIvQkgA4UJdVYcKum/U0Hk/egPFJjk
TMiy4+axYrlH9uiCuOQhgNC3loR72et2bTfmHrRIrfVGG3+blW48W15YADdIkaWOiy/gYCKpEcM/
xLVoEiFJZA3tnw5zWvhADpriOwR+aboj5CF2JV+ULlbM+290jVo8EgkdZA/IV+YFTRGJcAOXU5Zc
CY8gJFSgUA203jJm8k1u3oLUmpP2WbsW9UDMd46lKfLfFXfKzxV0kds8O31tln5AlXK6msYrp3AJ
p/RKbWJWVQoT9a/K+JvLELeKVGORaCF5B3ZVmr4u7eDPGsD6O6b6xiTkgIx/S4vWFuiwzswkNRaP
BEf/0SNhYA0DPfB7QdSeZyNtz6AcMJtB+dQxj0nH4K8XeSHfzd8ubrtAeV3d02nmlCnvMYZ8NPP1
J/VFQlsB1jNcdLOQ4XaWVnSIbtxIOT3HshKFJd4YUykrgbQp6LqcZAs9LFTD4GxgqJksyqPhw37w
vsZd75S/FOyHnvlTOX/s93yAmVXXfxLeVtK4KyxBXb47fDSdsi+zwMWeZmumDgmW8CfRwMngr333
77DCCeoQ1tHswtu+OO51b7moEg3ogL8EVxtxOHNlKcOt1RQKiFpTUXH+746JavPWvEKvK6KieWlI
ZjwP5zY2PS/2hL7xS0d22r4lVwGGLZtgIvc/SDAHrbmD/x+oXhzckOZoN7BJhYnLdU0GDV6ZCLx4
iVZzrS739JwVhuegrFRcxD6zWd05/rAHcGY9IV7TL72gj10dMxmhh5UHBNl8B7vlyoOTxZnRUIqf
MRyEKj1AYgfX0eAprx2avJpPvsXnrZn0IXgyC8pw19ogp8Bg6D1iSEK0xWgTmqkYUKnVTyVR1Usc
txiaqUvMdsh+aaMnVARS92n/x/x4xVhJ2eY5FYFXBseGeudrrFmwVkghyM+nAZKm0mARVZxnfdGW
/h+0JWM+VVpp5/GkM+Xwb2/rHwtNoHmwR9D+EFtDM9fjJMDO7SymnMTfNW2SKb7n8ZTvXlUp+pCm
MTw1y7eldeErN3ZZ9jRiMjfimgfPHVIKYE3MyHi5Pp6KyU5MGCt1UnuW1CqfiynFpC1VzKeqQaan
a39AfxWLaAhukWwvrpqZb4Uf8eXmHHHWLTkdJH2uKXpmxwBN2mmxR8Nod/bXJVanvWiS9hcKveeC
Mtf29h+HSHHxkrz3QJQ/9EvK7KaHlU/l1+HMGD1aDySgn1SlZS7+s1f4aYRNXcLyJm6YKXz8nAak
+qr5fv0mMQj0nNBPSwEmGUQet65tuyBsRqp+NY0ijvvhg6+3LmknGxVewWRqyMRyD8gbLtd/q2bl
0ZDmfXAwVUXAsgAI8k41dHpCawLHLuxBW7p6gLJsaaLBIGso6W4PrFHMmiaHCpROgKhtv7QK6wCR
2kwemn6sF1MpFutu4CFQ0ARsgk4NHUWcKdN8Me9zkAgpebrek9vXu8nT3IIKujGc7OL9w1xzmGXY
tTHkUHeNDLgtDN3idZ7fE+VQ+vnOak9Agsh1frEJr+GCqSYDAriEOQkMNCESWFg/UJ4UCkj1OsYE
D+xEAuf7oj+f+iXeHDel/QH7gtKG/vk3PXY9/hUgt/kpmLtDDY72t9tWBE92J/0gEX/UdIkZ8A/D
GizK7LCPQPrNUEnjwYt7+2z240tOfafwUmva4uj6KmQbotK6i9lkh1/S7ReufZWX7RfrMKSbHQ60
/K28HsDmwRD7YTN5jkTTGXWUMp0rkR+LKKaSNTeaR9Y52nEFP2Kj6PgnKPm3bhjLquSzihyuWpUw
BEm1s52jxN5Dk0iozvmrni7tY/vvkBfa331zxBm1h8GAqg7M/ppEwpK/oZPHByHL8jn3cqcAVM9r
Nj+yKKE369wMuGsWviNkOMkW5j4kNUUjVl70vwEsj/NldNB/zbqlLt68IZ7xjQkw2IOG9gtuk3/z
EgjG0+wwIKPDSiu1ToxBLjLKNOyb4f3xvNKL7MfDslygDOVXFHgdsgYUC93vEtGtHxjJL+doJ/s5
239GiSk6mYSodHgQg7GIaD2t8GNCm5uLwpyxr/hGRhXm6Qp6luaAqb6RP6mSuTfxU0mvTwOW0VI1
h+/7MATwhrYtXQr9G122zmldqWo1Trmuh1EjhX40iwIsuThS3cpD/ChkmsxdP2Rm8yTBg75CwT6S
tjzM0YZp2Zc2HhBloSJinHwQ4VvkUhfCv4Jry4VGtHAPLdZrpRC5/tydwRKY3p5BENXrbBadDA3r
eZnKFliYHswbd68m/IxHJvTKmupxFl1VFuunXkr3rvCXB75tZ3mHV/IziYVCyO7rJ73k+JgJWlQW
21uSklnmhfvs3X4iYaVxfp/k1t+z6gWmvue7x6UbKFGdkg6/GEsGfvPC3OrgVCN8pkHlm+KXgNlt
MDRkYaBMzQ9N0QAR5szRl7yWZnmfmqU8s29mNwlk1skjNqIYAmrfF6wg0mYdun9/4HvEit02EfR7
/iKOW3jVYxTRg7df0i3a1KxOd5aQid6HDwZnNqyj3Ao9U9VNiO2eQss1UN4OiJT0rjIkkWs0T9tL
WGXbU3TUjjC6NkDUHnD71LfOzET2ymKENYE7v87OzQTzPhX9bAVYcWNg0+eeeSH1OLju/zsoKDT1
cEr9aEV5m3PsmxRsj+UzH82h6B7zdZW5Mq1IGxUMIjRkWolvaAz/Vqj2mXAgbo+7giDRKwy4l8T3
tBpDaitqfwCqqitCIAkzBjmAvWzTBZlgdkH8afjV3wItVqGKCcNv08b6+OOLuQfl+G+j0l0RGnTJ
aQ8zapv2QHx5aKDzxOiNFCunTH+tcQRbPgPBPfvhP9Ku/M8SZYHNZnL1p58xkPQnXwupbYUPLa31
yXX9KlwI/HRu8hvoMqCL9wh63FvVoU37tNIzjjpZWokgzHZOGuElvsUPXQ2vkEUqy+ylHSxQk4TN
xbzUtVvDyBhSsuteDs2gorwpkV8CPFd0I83TK1wSRx+Q62+dEi1FnmoJzu1WORONUaCt0iABNFTL
l2waS41OD7uEJdpqEDh29e08PaFotJq1UTM84htANesyqaWi2qKPiJKPlk251eeFO25H+ayjeWcq
l2pWVStZun4c2PkkAER1vhwNUPQTSzrY7Sf6rbH34rvIoS1259KQVs8Q4SXB4hbq4o3fu4GkrONW
yK2d+PaAVdNMW57UHbmWpUzDhI24tGesVndIhmf4Li0/BRHV57kNMY+M5k8XdR9bUtulizrncpWo
qQU+spHDYUC+8k78tn+LuOJVA5BF7/bRgrW+pXlHif0q774N41Fd/rc/CHTiwZ9oNYzlaH1uCQbD
WGcmtPpg5RtRGQnUpVZCDlfK3l1zq6l0UUU67phfjJrbhKXRtm6rY97JySVIq5D28HuvXy9W9WF3
2IRfPXIZq0LZcDR2bB9bEqBqohNBxGvawwrtR35Lq6OWAcoHAuPSMJgP2D002gqAgp/7aILgX3Be
uS5ShI2/y7Dma1863tgI7MNZsmdLG9bWZAPE7VahborSu7KERHsnkGIhLMcl/fs37hTp1TtmK4jo
NBSpxK3IRaSN9sltmI04ar4TFVTaob70gj4Aer4LSXcrTN8VNfNqDvK0Y1q6a8ehGoN0Grvz84AM
AOwNSwCoIVNcZz+q1dYnn0+KJxzal+KORiqVZSrJ6bVYN4+9Nt6fRnoaLlBZS+3PFvTx9ije6OcR
x9OnuHbXpw080MUivexr6LNl7ZsFmUhZwBJe/J92SKV2AovzxNXVVIlILJ7kP5IG0iJBrLsxQHW0
DWqTlcgknHumYddij2e+eGzdWjJAk6EgJCYNnF/DRsKhDIgSmH3ZXywWmnVdkcwq47ZLvtsaX6ML
oejDfuo0/AbNnXtrejxgowEU31/DTou7/74957djgY3sPuFVNbs5fdk8d1qWRQ6A8je8yoWsfNMW
X0ziDlqmd2LpQkfjbLjMcv2A8/kBbuqsStIx1iKp3BW+8w86cVV7BSjYp/x7rsG2BtoHC3HMOFvi
tt2Qrzzp4H6MnwUvMJYUBzPoLwFU9IMB7QESVL4oxgvAqAFCwn1nsGcgPjC4ZVr4fNdHaHCNB5Qm
4B6KIGNbZJ9uKungv2QeDA9aaCCAOBb1ePlDdNpOa1IIpdBjwIbsqNOc5SksOcuCuxWCwYMh752H
sM0DWAezjLiZmZZXuC3VSs46xf0419AXr41a3AjyGizXnKdh3nfj2u7X9Er1msq3UZFAO/FJ7+5J
yV3EbJzaJrZdmWDHBWMAmHp2UOtzYCE780GVJv99XoO6laVJYhlZacOULmiyPI6aMztf4EuQfrIV
q3ejjtmwYVMsBjlM/GUMTOgBcSF4pns6QXUFwjWN25dtrXp8ovBBam3GlNw0JUlAvPMeMpZOxww3
rOwCiSYkRQQLSaxvdmpRKr30qB5qKjZjPtJGOJNcLCt2M91y0Hu6Jzbkefe5sDx+/ajLuV/k7aX7
I0La6r+9WyAJAraDsdk85USP8pRNuFVuZvlE1772STEnsZdAuCVc0A8tqTwXaTJEFqcMWiVCsPT4
vGejMxiGGvJh98sFJUpDZgzfc6qtJ9lnS0m0yLQ4TMuG55RRtqG5mFk2cwC914dJE4fExGecVQ6w
tJlTJuhOVJmCYJrs3Ivb/4su/B8Vrsyd7Nrm1uLwCdoGPhh+uSVkgFZCJKZcwAcRd1wbDXV2Dpfe
5NF/lGom+ymNrH+6WRaFtSftc/XVobaWp0lilHPRvM4/0ayscvxX6IyjejdBely9M87zFZplQlqw
OTI5Y2+BWlhzkOa3HO1Cazjxqvjgt/UZGoZRA/dm5zu47qL14aE4l04oIF3tiqF6ersoMTdDyJ8z
JdKRkRjUYeMgjAVnT2OedqLSBNJQtBc9QPfWdQYrURVgotrjY+pM3Dd2A6E7tDSJ1DuJpPEq+qEn
YLzFBf/qMFcK1wd8Yt/fRn0/4XjKXh9mWmGvltPtcG2c/fbnxRnM8DQAw4nF5MBL/PcLSU4ayXtt
N/A0sykPCACUWoCl7yMc8qaoMJ3R26CsY52/YpxbEiav0pPHhyFmcVK78Cm5+YASivY2V1UQeguH
aBkw5aJF+I9ErwVo6uBWXGHvFK+CTconP3K7rak0yphoxEtARFK7a3GXSgXBk8GnX96MtoxBT5Gm
pK3DoReaqJWGuTAsxk3oE0EDQr93U1N22fvjfmaEhZBurydkpDiUyfFYP7xx06dILCqsmBqYaX3u
1h4oFpIm+93sy1AG229AhbWVrSbHnGJs9VAAg8FvhEluiPjdMqJ32NPSNMNoSymNuYzpuOSS5zkQ
68+QXvV1G86YlipC+WND9o3FQbQWUtPTnLuj0Yc6NuATEbSzPNLneY/2F7Xe/5Ohy15Ad/EqXYzu
MQ7G3ghTvHVnx7i9Gp44c7+cM+yRm8gF+Rr6hPry5edaL02mqFIYRAaWYLNasUwmIMLyTb0EsUgO
OlXSje51VquoiEEoaIPj0tR2dpPrYcO5J0oiEbtPxA5SbEllx52DdKJMEPcoWZoEwItgQrpDmrLJ
0RkjD3S2WgDqyHZ5dwVEUDqP/uU3AgVAHvSyJVLx4/+Y90oLVt2mUYlzNisuAboSp1IIKY9hHRyk
KuNP0BYNuc3s3ncDRpi27qFP4lVW5SoZDvtTw8s9RjMsCxfNoChcGy+Naa9WgAWufUTyJweZR9Mq
TRngObP0yDs0E6Ix3v0aPDVE7EIm4ASMn3WGv9g2NXal+mSY5hV5AhaABCbou+dZYC5jqrZQ1mv2
GTOEfN0WJDN2n1HyukNZT7HpUReberz626Vmt2Z3BnSfhOhiI22zIt3TDT/QrI2E40Zhr+RDb9sm
igLhWqqeuoio6HVB9pctporknhZi3fj9DdVww5sh3KQVsBWiD1DrgzQ8zvXidPrSWRhsoX0JTLzO
49uFBlqu7o3FI5BBhyLwPx80trZGID6Duf8kXQLBozBJKrAYH97XtiFq8/u41Q+a+WhsViByqorY
25Tn0P20bFpF2UkyRcr+Z5nNTAgB19F0cLI/56GihSvB+yK0xZIrl0puN+uEO10m0seLdkh2IemC
nL8BXl4DCHPM5Gx6MIV4YOuax66r2aix8ldrc7TGwtiG+swbZbu58krrSZggzFuB7gUS7tANq0KN
BoaQSJiOofzFD6RlnD7QpJazUzRg7tX4dzCUpt2EEfBUDtAiELdyOrLIZ00XYeqReUtPjFKcl7/p
OV179XcWQUOYM3R4506HGxemUr8/NNOrdzlvqT3FT0jG5tDVTkF7z98UG+ZJ2NuaceKV2Z45jhju
vk+AisBX3CBFFRy+SPMfyLT0tpSmqVJCBaoJTLdylHhbiNtmvKc2pbXHr+c2Fzr02AyJPBumeWtE
nlNnlrw4/L8W8Ku68U78nn+7YLsJWC1LZWxmOxQ5DOZPD14f/kvXwo6/Je2qTTUs8IrNjTloGTF3
jGSs8didbOh8oFChcJ48hDGuALoQLoJhxa+1D09O4tiFb8eFL8ou1awbBHm6hqeQ85/00AS2qOeO
IJVUXDuXOm+3prjkqyy31NrinhuE+g2ITsXxjlXoMfXAfMfqcCDIojt5Y5IoqcPQ85hsSTA+KoIG
XHGoFGz+LmwzrHNuHqRny0z2EP9gFZbJn2GkyJdHdJt8WGotgC/mL+LLf8TwGIY4EO+MAUe9msmh
KRMjnlZLFeiI9iK3JV11muAbQkMvjfDQ4h9x3brWVuleu5w37Vjh5NHBYCyPKSS7H+VblLzTU+xH
ubcJVVJY8VCyTzYDrd4jR+/eD6FeFF2fNnFty4Sb1dnQUr/PKc2htm9FCJU/LR8HBsXUaSaZazwj
ahwHQi26hzgYse1+o3hQN2yHO3mHHQmr+vhisM61gab0lcy831vOisqHT2uwVT0MRQH9nuTL+mer
+kBVHl4+86ptEHh9UrcfGjhsIBsXzAnBhl8ZcXdy87UO+k23R9igc6V0R43Gft/ZFKvby+xC1bqR
xacCFTUC8bVMPBMau1NVOvusKqs8ajyBw2s8uLAIVxc5caCKGiIR+BfRUtCG06tXDL1FsSpitotm
5BEnE5Pfuoo1I8iRW4tIjWeOKbKtymuU4OWnF4/9tpnObW6ijBrog3Gby8Frz+opIJ5ZuB3HIquD
LdOgqgV/bYDWBaAiCrFXPysSWk1WK+Ader4mwsz6Z6S7T+hEashtLzUAwSdMTGEHxCaOEB/LENsh
8deDhmxoBP2MuR8Ub3cKyC3dIA3rUyYGHDSVRF1qLSSr3FXmlG3Z+mK8e3Fgm6KO+KYg57i6hlZB
Ds5dwo35UvfFlhXQpv6GZjQAPy+5V4cyQtaEzp5zmMUan/cendoOTtQpsRhU+0wW7lOfT7yse1nx
Av3k8tijNmMYyXiq859hkHxiOQVvWdxQdh3PYU/rJqHU7IxEt3mR1BX04h6RNLYEMEVi6ZQTQjCn
wGmNiw9RMAjd/uBajB3Fhz/mrjwonv9gdaRBAs4C8UCzv0t4T+uSo2/6noKPrt/nsrMW/MxbCNIG
bsIQRyjz92ImZqHiDnWyamTJ5rmQfh33MKc+zdpCzdNJ9hunk7ZZupZcPbtFSUs49EyS3kp+bo8A
sA3pmbgzi4x6myjQt1r4h+SRILBBAI2rU+zdBlx7NKeQM5rpnjLKWDxIOi1PKhv1BIbaL96DC972
DUep90cStDZCHDOqsUsoyH7hEOCqhJHrIIbOainwXUrWgRz7YIzLls9SIObDwBKXuNmh68HpCXMf
2j383LiA5aqhp92mTKC3vPVGAuvrjwkzyECk+7brRCQFwdwE2dlCsTznjbqGBPKzuZnSnGBxZGUL
nS/8m94kScgh4wXTXo17aul7JcEWY/ARBcjdvzS+PHsUy2rG50jUCRXOyXmvcfUy5F/ITpC3zKCw
P6M+gAHzLj5qZeEri9eJUg5xIXC4vlSxYGeRGbSX7kMfXNvqbTrh/jy+KYfZ6pyxT7hbz29uoM2C
hz+6i8VbfR6mgKjfd0oXW4PybTtAR49mrJ5GbVQzjGCkrWh1X77397Cwf9p5ecE8uvR9nrZIZcwd
5rT1fxWgw8sTyR+xcpSokLrygeSjO/aORIV4I45ELSEsh5qR3eOnKfR7x6q6o+UO2dbOC8oqFLh4
96Up1i/GlbFvYz0x4p9fAg/GbK6wEIYE9Yv6lFakSzsm8QcamjCqchS3hRZNyPMXTTMEtLVutCfm
bHTwPrUQctnKaeMoBFYzX0qvS6r//tyTW5OpET4w9rqmja5Zsz/T+CzjfWS7U9ya7B0d2LnW42kc
j0hwDOZUd18bcTGFqdz39IV1zjkk0kyqAmZ2qqlVemrPeVWgLmOnybPJ0IKeyg4l8HD8O7Zn4eU1
/g2MIKyCuiU7ZKLBcNccM7YACbpFNnQgPH9ZplnrxRoA0IpPpnvr3NNoLaF4t017vNfeXZ5ypaNO
5kZLXMvje4YYEdqo0V8059xVq4B+RCetCtW5l+LD5suV+iK2Ey52Xty1CK/R2IzWo6f2UMMgUlrX
9ap7pat2X8hVt1BW/VDfJEk4jE9mQVOWPK3mjAJtBiiCIjieWWMKKlw3xG7E0pbh0tPFMquvlbBZ
8wYDLV6iLV3CHiOJyE2JdgJ6vIQ4Ov98MpQ53tVEca7Ob9eok6SgL2/zUEUVCqBUCJ7ldjgbUlax
7ATB/C51ywnUO5oN84NuSU8ANcrghDqFZONMJlFg7rsAESSHZnHagxWP3gGdZ6Jn3Pb0sQtfFZej
egGtUtgfbH6dtp2TWJuzaiFFTRy7joeyTHHds2wfNGXVu64SKH4Oh3UrXPw0pMEY9aQ9kso+NY32
X4WuQveUgfgfvzPNAIA0VcmdpJAl8OSKLcXwKDkWwdXSrOtCMOxF+XxD1vPdxqklS70YPfRxap5W
Nc31To4oVV/EegYNs2SO+zCLxq9q8/+XCRIxb7fqqduBXPRQQcuV55YUsQOVmsO2VdItM/GHqTTn
rqEtKRdwCtBFZ6JgNMMOrj9m/HpZPV3QjnlGbm/9MfyTEJ6MCHXpe9ddrgN2p206qdVwz+yNP33G
y6ftsQJ2pmQjPWzqO/QsCc6XjtdCSbl/3jL/o+2cVBPcbjG1/3vdcYZd8NeS5+O8UuNkC0Xj4AlY
6CQRJV5AN9Q4skOz3IO+zPbVXO3UoDOrtVEqEBlYzMvPIu/fYTcwVdgUwMIrfIiz++0ZsJ2z0ZuC
Oo9sKRXpChyfQ2dIb1qNYvZ1W8Ufxg3Zt9dxt68A1jHCGCcTLgJ8wkF23SwJTXnx4qh6eQYfwE91
IwJBLma5FHTgDSCEa25u9jdsDAR/qFx3FKkaCIr3b2FvOfITtqa0WanAqhOfPIkqiM6YQyqi4/hQ
TtBUpH8ilpXwMLAThWS1vtLoKmuxwDYOWPgnG95A49TS78tbsKVjqDBQiNfTCUsDH2LXqMnlfh+c
LCAMINFJMxa3bW9ebIBd4BoaOxJYgEubj3K5r3Ezt4p25BYGH6BmwH8D7iQt5fgubKy82UZTIWUB
kWRu35tOzPqnAwqe3emTVnQWVTz70VJZtFFHKyuGsL6NwDkSnN3e5uEJ/usimiySqKuLzysrql7U
rfHvKS+hLgRenVp97waou1ig7whGh/XCrKTtSAHWPX9O+r0uYvSwimGd5jzkYkYxZkAK2t3EmZQ3
CpjHbM6G/9NJdqP7vmr8a+x2auzmjfSSgtLANGwduwzFE9Fb9J/bTx8uvpRGFOlfq3RBkR2AgFDy
Jq6NR85rgk6NH+ol+0rX7BotG+VEzXj2qAgz733t8+Cj6o/68YeGjG4KiWxpRWeEarVQAcIV1Dh1
+QrMA85wKmi/aT3uf0YrkBHt7il2W1uyq67bj/TR2Ax7SkletLKC+RTA4xpVkAHx2b8QGJC5dMO/
SP4Ut+UMms8w8TAlm5bmf7TrUxUOKBQzhbF4/r//d30BZV3fWwXg+AqaOarAxLl83uhQ5rl+qxDx
jxcRXgel3oBSXr/DeSpNArZOIsahnQQe012J6mgk5f2Tp2HBhSIprj/hzUwAqVB3v4a30BqTa1fv
rE/PGr8I+2W0p66gETlLD+i8q6oxmCivSj1OHG34TrY3KvaMrs4tIpmJq5htl2rGVrtd4wA2PrJx
NvCHIX6jpJy9ehdavnW29HioB4OGGSs86iGobXEb2YbKjofbV/pYnzXC61Y3MnMbHDZiRbgrBQe3
T9hZpGN+C6GmBhcGAy9WjbRP7tQE4TacJvDAIRx+ffRkTmXlby5iABADRc6UXaG9eLNGEHSG4l8f
Jz+vZb9u68999r10m5+9toiPJtDNCnQUnm+krljwQyaaKaQf34oqe/1bIFYNYCtuO9zq5jPBpTFz
LUdUxGsDZGXFCNUU5/PbJzSaH2+gkgR/AJLbf4NhInbHrnFf80fDT7uC+zm0yWhuS16djlJ5H5TN
nlNrIk+vT3bezpfpp3D2NA94kAZwMIhybiJrXyJ8do+ME9ZfmAUNLYxi4cmJVzx+s1ks1BAPRSWE
f6ek74ptLVONjp+QtzZRCOFD91SXVuNMe3rp36d9QjeFO3Orb2GlTk3L85b0HZqQz7CUkEZymZRj
Dl2ohrF4EGVx/euPod574VneStGgF+bJDADUcECnLpeZcoPUdOfR47q8lIAXoQvQfCzi6b86p2Pq
1RaYlq8sduS2etCfK9ZqodTIIg7xRIFra6vQ0VOco+Ox2AwmkM7F197QUKE5K/zMOXtNQwredpqj
9/JmHu5wtMwnV1maahxY0z+Gen6MC+rmdmmzlpnkaW+N0rqFI3pvHaS4HHij466tTPNlyvYTRR1+
aI0gLfl7S1dPQH6Pumo2dLuhfClu7sqXD2DhU+1/FxhI9+RKi+LD1ca/Vqx6hrqyrnIzKSoy+HvJ
tHS8I5QSVq10KKWPYu9rgjVoPVwW4gIwG1EPrJlu4F+x36r+CwK61TL0QU5s4jTIg0yQSMyo42c4
WreWJjW/llJMoEQKOVuhm1LTN/Cpx2D3g3H285eMnBYu4n07c2ud2FsbfS1zepZRJ0ST4JF8zdcF
zAyiXEcHpRDVE3Lg+Jle7CPD8hXXoDiJjYVGXs9+12etKa80jU/u9ojd1mFhrTNWUKtZLZHvGPcJ
2q0gc59vCpkJrSHkKGTMMMs8peIAeIwQEll8XVQ77+WIJx34k8DrzO1fXC9PVUKqvv9mT3wvQUuI
1lWcYDxNixMd5qKQo/LY6dgNVgrSibkgiey9tqQIyoFO3Bfy3gAxNOTXjDYmkFQThgmJMWhbaEvL
GgfYC0q/xybaHrhEr5Qu10+KL0o08V5Gkb8kYVBdkFQqrix98qTikydJAA3dJ7zyGM/sRR8TDl3N
Ls4A9dxzMPkuJy7CLQ8M2KHiCLj2mtjZ8ECxWz7MlACxxCKcQP7pEmdJQ2JpHEJsM82lYBZ+9Dze
iPjowV88OWa6yqBFG2i9XlYJ+1IZ0bAn1Nzm8TQ3vIEJgHOTHF1AcGJnEKDhlXehjwwe5gFebaa2
HEdnj6ibXzvmDcn1hSmj5aLjKsPfwGWS7hPANexezjaUwj5VwctsR+GDlES1MYxjEZ5tSObKsMow
uJhZl9zEHsaIFZ/WBDBbDgyVwSLTktOB3Ce2fiZwGv7kVAUBxPlI9ACuhm1f0ZYhg9Iq0QOFXou6
0QRc/vQVUVzHNdYg8DA7lDuaumEi7KpOOqKJ2r0qiU9UBEQOMyfQxeAS3KB20SIVxNy53BoyYDZT
pg4CNs1FNyRKwqGCKpe4xlE2V5up5JhqkzUvqriqC1zfBWO/H422vGD6hUFp+sVIrTdNDnk4NMR0
PCW1x90tqkLKQhjPwbpzHR67xeP4anUj3ye53BQmiyUM2bvlngImAY7/UgzspBAsnvW3MBHhPr1F
dt8NccAlJmwM82r4mQAHL318j1feW8lFypAZi1tqE58KNLyD1BRj4qtLkR4OUqKlP9gSKAHi6t9x
d4zQVgxVGe1UMgSFS7XKkVCmxIRv55qTsypLQHlaR2Qc1220T2j5rv2CQshqhfMBkpDj9MeL71ba
UuYfPvj/T8NZB+BhJTcaJL1flspmAY+Nqh115uQttCuMkWieCAjmmAfw9qrHlvntXNh6Tdm0tZW4
JiIzdM0ZgNOTJTu/Lw7Rf6T3l6jqdy7Coy+4Z3Wb3t6g/5842oAT95bIBEyrwTMmXArBv6KDdgCh
uU778XnFVvqT1Et3kJR1XWBrhQeTBOeBnjWRI98KOz6tl7Dxk0zjjeAiq0fN2L6Um6A7LhOMXLak
86BueV67gaeQZquzQL0W2Q0UTU/A/+jDOgEYjJOjfBXWjnm/68QLfVGoqvS+zQuQcrHHVCEvlspl
IqrgFpDNR/YGF6fbZevH/BXB+lVNEy/NoDHdezEBuUfNzT0SZPfY2LWBUE53JURLUXyqasipywHb
xRYEEsM3H5N1qUvEM84kaZmBPNjMFt1XK94f3VVfXeSSt4o6S0RhL+cUIcDhCV7IbRadxch5Zkv/
hOMKRWcjSZwHolsKDCoY7BDFFfWHoFluoEe4kI/k0fkJgjTpGLN9VEWlvX86QDHVxDy4RXsf5Xjl
zDGtVYmedEIewpQZfVLNB5e2rbay8LqrojD0RECXImicknuSG9Fe4SCVwf4IoLeKe4nCk5Ojr3hA
lntcKDSgYvFLOAxnELh7KL53j9BjQzpLYbwWQ8On9tCjI21/AJGTjsX4OJ32n8HzphBF08lvXfO8
easbYXwyPCdGOHNltVrKmoUxXLH5HC0Gmp/9fgyCeHxFuILHQy+jZRG/cV6eICZr7MhJQW3qtxmg
yx1+7o742foW6dNUfNYY44TTBU3JoIu8kNMOr4XJ/XeUeV0ddX51pM7PYaOlO7RbE15lb/NOmYiB
TIbQqWqGNuX/khmEd/YKaj0sZKFH7ekD5+xiy/5u32KhtefLCyEqvAj/YE6L/5Cg484eh0mIm7CB
UFc1N0mxSciL+qh79hPrIYMJ07TW64G6g6ut57Xqbh982f54t9Cxy0QA4Sy3VoBQhUxtRP1Wbk5/
hdN7IS6fYPlNjzs669vcFtwom0wjEkzJJfEY8YobZz4cE/9PjtLJ14yZ9R5WAAwNO6BgFXuR9fFz
sYHpTB61TXbveQSu5wUyaujyQ+6nScIy0GPVNbX1hSJ5UnHp9MAaBTypc3yHIEXjAmiSs44TnqiE
6dHkgo99Q8ZN+jXezi4W1pUQoZ23a38ShyeHvfMRPeYAUh59+RbCQNk4aKxp2obGb2MQYYGowSVw
Nc9bI3u31IUEMRqfuBbiKhFpCeKoyPEKinsQ7WZW4YFm06SGm9xHbiW/KSMu/NlZHE8rrnYbFT4f
/uTR914yu+ZIt0dRiEUItpBRsYB0BLrctJ8jMVfOS3e1gWSjNJh5JI0I668R2MXCWjt4Mu+FfSON
3B/X2yzcz5HcpYbVl6EwEZXrOxzU2alL97MRSV4Tmrz0M5YdvyAZjSCCRX4hsoNnBs+EfmAgyxOB
zyfwCn8fckjHZD/vQQPclbEE4YgG5t5XYajaCpDI+ZW4+wgDUg7qIJYdEidOP02D+7PC4P6t09Iu
124FfVugb/fzPDFbz5s86rEBdaY+iHbe8w+i8E8kHkQpD/Ma34RvTbHheS9qs6HXVYbCqhhkRvrY
Bcs8HFKFxX1Ge8F01T6qNu/Ut3b00DjvawNhHKFygKISf/PRXFPdsBF8/4gta+m27q4pgvQUwHnp
yblRnYpfSQUSHew+xamChd/q9SXNFFsIPi7tZMdidJ1PmoXjeCQ3r8UhulWWB2VNAspeRAOgVToz
dffuy667C+T8SckPuv99xx6NB8CgTD0zdxGucZ7dTgXDKUj9trTklFGKP6XEmW2VHuU9rDhjM2hn
kNDTqZSgQ/c0CJ3LsRqSWmmOoIpuByuvr1rYFRzIHfv9+qb8WXPfXXhdMOeSxgjfe3Cdknqbb0bl
ItGzTJMVMNP3+vP0EAnPlRJ4NG3Px2f5FnOh3fglo4HrMf0OkcH2I41ssGXDxzbjhdPSG5mOq4tc
zjsuZ94NjTqY9LGUUsf62EKf2kypa0mKRHfWYON9P17EJ6250kPRui1BDrBh/EdimjGznd72Imnz
iTeHWUbr2WGbsvf4HHmRMwYbT8GQ/YwOXOiCPwX7Q/ub75JzkLYuW1iroQ1h3krfujhR0yvK5mCt
adYFKNzafqffEpjDE1uznldAHIlji9T5MR264om3V7hXuCY0jlcie+E8nBozjioTXM4f8u5/GiOD
LKFlg6Fy60kuwPelqjCW2pbiTfOcURnZJnmqWlpMrHrI5IPs0GiesDImb9iPtww2cJ1ozxc9pXZY
YVMmXP4NK3KdfD0VfaMMi7EPOgApSwdJ9ZLibIslEU9pNitdJjjXTxDGElGBoKfZ3RJ4JPp/YM8S
h8xfMOUzyzzHujqh9YcbzpgSPPB1kQu+Gn87dIj0GUyBemE51DrWnXbTIlUkLa1NYGQb7ifTDa7O
tN5uizfaj4MybOap3wGriIynMtRI0jNkILca+Oi9CuSb/6O1aGTzSZza6Y3s+Wf1RDQdh3G5JvfI
94kyBxHCjLo2hivvc87XXvPDMcERk3RpncHAVB/zu/iGg2QlzQWtAZidltBkAqdfM2GvfjAltQsG
rHl3jjWBGhfvy+1C+Zij1ls/9KqZVHAWDX8TWjcpLfhhJj+RVpGbDeWAP2jOFgHsWzDCwid6kvVR
4M8RGdE7QgWlBVr7hTSJvgUydHVQEZV/fgk2EYaC6nKDED9Jq9tG8WUl5mYSw76IgcrUbFW07dQT
7Bor+tzZxRtyxXKJQS3+q1aiS4aG++0mRggp5Gmy2qWLe9ka4URXE2kv2+5JGoft2l5lPWphtZCX
XXn62kbX2fI7kCMu5p9XNjR13WIDxIDE2bNRbjhxkoTVTDsqwWU6XpSap3zfc7/+R+uVGbnWuQdW
YmuwNpYJwaZZO/3VEvDWdE9oV/y3zfm2f7ui5UxNDycAJmmNfJjzD20bBpDyERoMuCoA/XMEY3y9
sgnVfBWuTAvCxmSLlHihXh+MmiKlRm1GQ3oxWvPKBjehOyyjYnFMBlRr0FKZt9YG/ioLsr6bhuMs
JmvWcpsR2c4u5fmjKzLLdmwgyHZZ2r99TQg31m52Q+3fdGikl1cx8QFqWL5wZCKxMfEl+vFQrOkU
J7MetzsFgB2IATad51ZXUADYqyBodp4sXgabvoHLrVorVBzlVjvy+GuVZCNJCXgCBs4oH3V5ms66
7RHZoDbmy1K7E7NeupxfaEfIBLKuo1JTrH9ti30MBdeBOf63O4lX2NNErc3KUpcfaPD+2G+dHEoI
G3tetCJgnR6UtbF38s7PzlI/m/0dWxW46exNxZ0ThghciN9MgmiBnSzhkBoiKlicHwrst1HsTqNW
rb5erMwqNOfMG0FcZGvz70EKzCmGmyHzpLat0todWXuv+VDY/IAhUeuNuYLPMv0kUUuDqjGrCqGr
XmngSh7yrg3tIf1izMBJtgLJ/6W+h03pf4QTsDxLLzdvinIHho5aum2wb61SCkQ6xX7u6LAilR1B
Ar0+5m+nguqRE5/eybyHV6X7Rn8NFKR3e/vWZBr/Wt8mk4rG3lT7HOwf/K4Tr9nuQAIte95jkiMx
4sd4Gf/q4yhV256XsybdqNPweHWj7AwVx3/jTt9EpZBKFzFdovHIflgZN9uMslNfJ+VZdKsnVSw+
hEGB/iZZql5fW0uT0MhDkL0w2y4EXEn/EVt/DSXXQOQAwoAxx5xeWvJvwfHZ60NiRgN9PwZPguqH
3IdXoAOHWdCnz8lxluEJ50auRU0WEM3ouO3DmWuJwnf5g+ebXx69bOlBZonnFnaaf7ZZcTDQIuP4
4E+jJipZbPaVDlFmZLW/pE1K5uMFAUKLgDcg7FLF2+twWBNMaknPR4nh2k1Bo9zxyytKVS1y69Qb
z7iXDTzSfibB5Jj8tUT5WlRgkUe5q67ppj2/gI98PnfaKTuK9gQdSVBySUWX7qyUwwdO6XkO4jgk
olSym6XN/bTCEcFja6UuxmrZwfl58SFeOBnMiUP9qPMgaRyenGA815DlZKCDx6JNBXNlGqQyUeqc
UX3Ug9SjxdPI/+NXxPg9CRJDHznH/UKjGyuUijO/RkqYWHS1gkxSmbOnJJsIJzUby9+WK/+CY9S/
qx0SHvUXJw4XhzO9A6Owady6htZ7CS805TFe4PCwciSWDE5ur+7i6qPr6x4GogYxK3wHQcikifxD
Sos3sx0S8IuQuGnL5aBIRzgIJnzOldPDdMqqoAPcO4m2Ewxt3ivOz8n/xxqyF/6re0CDmaQQoTD1
pUvShW6SZ5mPL8RMz3HtLsfajzeJKlr23g0zJ+xDnzzxLc8IE1ncO26UYkF0NMfS6qRllzOYb0qy
3byENd4mbcz+O8O+ASZS6FCY65RsBtPSvLN6LbSOpsJrmcDBNi7yO634W79Ao1Mvn9AGC75uDZ6Z
upetieQadsgF5riHwD5kaH72IWOuaJqqa7TbRi+u4xwjfZG28cZnTDoxjok4YvxjM1dx7XIgCV8E
JVQUGUXTnX0KYv8YaeksdGT0T3wdLS9kdnxV7pfbJL/mOpAZXrD1VQ+CKEe1QwW+j5f73oGrm7DT
1ThE+b2jOFN2H/AUlumUFfoalWVr+BoFLayxw+UFvEK0RP6SUFTn9g3OfJ6pI/3K3Zt+ny4NjKE+
z/7EaeXEKa/4s2tT7yFDS+lbUCv6vRCj/2sbAccmoqdqVdsqN4gFUCrhyN6OzZMI4+c+maGf/vu5
i128PukgSEaBo5/16i47m+fEj30P6N7gsbRbrPMUad5eqHvlz+8TwBrZKPQwxOgXT0y41Zk/sDqT
gQO9m2+nYpsO02JGTOdy4o9rL9kSwtn/WapXIx0PGGAxCRV8q1eZeitaqnlENGSmbChLm8Pk0aeA
N8uaiIrG2a1nEKvs23RC/AfoRPRi2K3uJ5DnjcNLxrRNE7YqbwiEzYGWZO2ohzQuhOEqMVt2GtTv
RnHmQDsLTzGsVOyVFrIXUwRTdP8KpgI4IlWuyG8oz+dAawWXAbYVGNhAIR7TpVyZ/Pqc2aFA9M+X
kZ11LoSkEXeRfr0D9obdq0RXVOgZK6ShUqWTdCmz4gJXHaJQDHynGYif32vPZyKcGHYOuZS8zOxK
99wyzgdVuNSvbnpnFV3twNl+0yBt2i1oirNCjNgQZ4BQEYsKs4s3j+GMljnsoRJzr+ydY1eZUCIh
c4n1sero1T+ap2YN8Kb5s0N+SRX4iHzaShg1OgxTPeIXajI9xF4T7kIqhPs9A6Ld6vLriomn8LgX
hFLZVXEfOKZdQaUch9ISYkrI5hV4bwv14IAmSalLg3cEqyVokeJzH/V+USvcljX35jXPD/jQN/+f
A2udI3znJ+vjFdVVgrbGGYDzU1LUtJn5BXz2hUxX5dzawJpzpBicJl4Uhv2H3Fw7uVxSa/lnm9aP
gg5azLiVjC0Xqtej94csxUQj1GkZhHINx4ggiLMByVGkFcLxtHCQvUie++Ujc3PpD8JcywMhn+/n
ok9TuzmcOlFEJxhnoszfoY2yZiddE6uQ9SRJW76u7X9PvsD2f2CUNRIFSz5WSf+T5egGqCyQ1EL/
Ge8YbjjXTWjOU2Nc7di+vV1LxpAhNsTAoD7zZ3FnaYAa7iZixAvjKaazLQmDyinbyNGOcshqQHD1
vrMKmapLzdxjgmCkAKLq9JksvkTP4RHpL0Tyzq659Gvz28bN6pvk2uf/DYi14glvmzHPf9iSO/z6
R0AyQE55iJ0JwdgINOaLN2Re6ja1QUoQ+6vSrAjwd2i6rGSDpQ4WrqfZ8wVxdAL9N1+A1QMrM48c
tDXaFvelPEK1Gq4S5oaFhaIZ5M1mc2PCRF8moXnIRKxtpflmEP6Ls7WewKpZczd/2KDDOmoLAt/7
9xjxQ8NPWRpNUuZs4yznAUm1U0wUQVi4VXo9RfP0w/kaLOk2Mnlh+uuyKwTLTdv07L0QUNdMsaxv
DKlvEqhMlZFNQgSlf4rJTkXfous52TEBXMB2ynK4/tk511p23MjG7S+g5kPVkIZI9EGiyeklgrFN
gK5NARH+T1hVw190cI+4so5uG6CWiptZWkmqJ9YIAB5Rq7YYHP0LWgvp58lx+k0BPg1JSOCTo6ua
cPgrpPO0/87g0vWnBlruN4LtVMd2aMl01aHMNQk0AMHGo48IvYJv0yMMpDwfMpUt4RsJ3cgvbR5x
ohgxSoCsYRSDlN1We5Yq1hnAkgao9hutTjrF8fOe62S8TSQq5dDMFQeS1zZJ5GXpvtIxcCP47lWg
DQu4/3Eeua8P1C/3btGY31vf9cjlcNquk83ejXpZRIJ0sn6lQ+Y6qHhfHccQbREfai6VIS6oagZD
y7Nv0YtHRYgM6D+G0MADtjfVPvwYZD9E6o93Btory2uZbgKce3BGcObLTTdNzjzkSDBWo3MEU80Q
euI78WGhF4arN355GwdyGIiGp6A7QOljeIEW+XwGKwb7/FsKVPBRRgV0n6eZXGRpKyClU1aAw3uf
fU+H700jwbdQ8wGJxTi+8/PZMJ9mqzsQVb4IhpwQWIF7YEsrClYiMPpD9E/la43PnQAWZrw5adqW
uwci+ZUybVAGlL1ynU1vOYF/kvWOGjN2U7U2IOO/MF9o7LxWiShVGyCc5vMPHGvAPiwyPLLKZ+SK
hPfc8KSFAGWjUKzs7Nikh3PLYH5/TsXO+RIBd7s/Jg6LVjBgPNzirLK/vHrJkyzfBSW8vg8PZOQR
Mrx13gl6sMdZpkMPZEBtOc/eqnu+HLXquovqcTihxUDKNktaXcxMMcwhqnCPEg5KN1sO2jY+OC5t
x1Xb4+aktmOkwn/i9TTOE0t6Z5NEuhMUotXFAknaDNMRVdkQE6MsNPqPUgKvRHXSryyezu9SxfVH
S8WJGSWWsHQ/oIc+7JFAkwu00QJiGr/zf5Z/Q83wFC68QElQhUjN2PAAb32P5ZmnggVrFJNx33dm
9Xz53GlwXGu/5wMd8pA8mFzlKibYSLxvqYUC9Kp2qOsOXcsHaiTSxnYJVqIfS8oKpcN64u8S2coY
thMMl3+FQ3EpB01xlPZR0h38qVagofv505da3Eo/yKtZKEayPh150YrrcaS7iIWWaCnClsW6eYDi
5co9xtUUjeNPkyOwT6NJGJ/yf0iWrVprrgn7M3uzNCptR21jPS3h3xvpQAjRkB4WTiSryGllOkf4
xucqngCFuAAfv5mAfFxVvF6XscwYKlZiUHYpSzm+iqdvXadgBCETheMbv/ZGOuWoV++t0YWEPs8k
RI1cbHXk5/iJ8gvOY5MxVinJ9fVvvm6/hgKXljs/H81GcblZ5b++wch+76D+Uig4lFkCokVK67yH
avkr9VLRQrT2VfAb9F2Fx47dDtY9j8xqdN46w3bi0Y51B6UotEbTtOQEkM9JEUK9ocMDVIYcK3T4
HzZCADl2C5S3d3p9X/lYc/oXNer3L+gMNZBsG2lhPK3OQsV5YOUp682ZpjE24ySU3L9Ay2kN6Xm5
7mqlRbSG1rr87sLvWx2a9rHklBjNb4TgClgExWmsmxJSoTFrIirPLMwfr6dwPk3TT/ey2TjL1zoH
gDEsc8nJfRl0hBe3tEcrLgioFZyh2cj0DUrgqnlxYmciBJIJyMTFqE2uvofAa37/n2TlwAKwGRYR
uFWrCtzo/vPSwyy65WjuFCVIwQ4OV2hOn6mZHjPzywIZRIko5avoS2n9bahd1x/wi8WXih258YC+
ZlbK5K3seBqhjn3YzunYHXKRYMGYAS1ztd7EU0PU0lHDjdZqoSoXcJYP5cGip5mQ8zb1mmfLofFT
cOqEVhwBiyIh/ZZT8IxJ4U83O+kGAMYIP4wcVLsUPKCbvRUwWPt5IFr6DbZnZDREVy2b4KZbT4uS
dwGPgho7mpnSDtAb4Uc9FKjaNvctlYHYjVe/QdQF12v+G1aVWzturBedcoNqvUj0MGoOZGjfQD5n
rl2wglFqNbUYlZYN8tqDdYAeepDumJUJdtnzu8HtOoDV3TjKxG/3uwz/WNo4j40eweV5cvyMkugT
7hlg2XNsPwrbuNGPcXAYabuuj/w736h0D/rR2vdJatCTONnba9HvOCqhvxBExwEn2pvGbLvg4MTP
o3K+APpklk4qsRgkVpar4ECXEjMlB0E1yv/pbN1vd042McBmyhjTinVTLIElHc0xPrlBnVnrFC3K
3zloH9ZqgQdJYh28fhtHMEkbdzzYvLaWzqPXUdKVGxk+Wvbjj5Usw68JEQ1ChF0W+5feGvAOnPW9
VcLqex8jJs4GgsZu6VUjA4u+YQvywAOihkYX4jRdy3wrKv6rN84CrOGM8sQT+B/TqNuVc5RgUEZH
/+RuilR6JjHq+Cp/oNzZYre0oEZbQKORO82s30IKQpK7uttZh08K+g1fWp40kSKGvgmt2fkf/Boz
bjiGhv6i/kG5X5cayuerb/u+avoTfPD/hJfnCx/HcUyFOZyq4yLWbJgwvSdc5UQrr66E5CEMRkZw
oSee6mx66PdiUZnDQEO6DVFpjMCqv9zxUnXe9FGILK4dIbFC58/nNCbd0YgQ7O7cmWD2sswKMXYu
XFY0x+MymudNOWsnENpQEksa6pYSRFfjH6DiIBnBW19rr+vdYr89cEEZ5LpQcyDMlfPw5NMlXrne
N9mrpuLwTQmVtTyt4ESEcnkSon+B9pCUUya2FX6qhT79fHC3jwWL4OpGlJSWPzkQdZTMjWGn1MNh
MiFx2uqamEE4crMqMap8kE2uidtdf60BIqRSNCIfZAb33fhbdrImlOeVVOgjvF7GBKViGfimVUQ1
xpkDNrmvA0pvfUUTpyij5kHaQvjIzwaxRcLTdAorbzTH9qQQw5zkb8jsL0bnkK2E7w8auQXDq1T3
Jx9WYJ7VbG2XBpjDEnhG7lmqJ3Q8iqAEB2ySPRcLZaEvuZbq0B0EkdLZwD9MYoWmrQNI3Yy3XHEg
8tZ9Jd45HF4z/Kjs/+KTk+WRzKdZk7lsAHbe9VvdBnIUSnsYxokQO01qWy5WCDV1JPqR+gAaf0vd
c1wWxd+cwVegkaAPB/LTZYsykKnoPLgFhgynMmS8+jKhz87j8Q+GKaEwjdJuy6izFMpoAJ0NGmzL
LmDLAvAeZVdQE2JvyuggO4xI7phCbH9oFWLAcodLcZujuSZgdwgN1dHQKoZErszzwqlH3hm7binF
6cTYNwcGsNUQM9rHEOOD0yaq46SfCgRhburxP9LS2lPqOM3nzQalzD7aMly4ZJBbJw828gqG7ALz
m8oT3xeTXRcnpHagLOimGn0CLgA5lnyh9gUCHKLnMxmNSM5kbNRSdwVGKqQtpz31/rABjagtYC9f
j/TpG9j/Lw3WItXIMLauof2PRZIzwWYG05pxSQp8wIeLJL0Ze/nIz4TqnZVfawZE9zORGOgu47PW
o1zkcGAu/hCzXm2C9l4Daxn3qC6OdYNDKpNcZDKa2WYA02q/S7/nHrbksLDh4tVkg9jrRFCeF2AR
tPsGm6i1BhXVCkI795r/2YKagnMoIYG7LrkpBrXg5LNT7+jXksV5FEOfj3cwqfMpj6OSObscxtoJ
xjk+QPnooAYdyD2V2PvKQa0AoWHtSsZb8+1stdMlNmFFfvwljXMTXhSfTF63VvqKBB5gizuqS7tT
UgI0ljgCNMlUly9CTGTfNX8spvKQ6v+WGnYepDy9+uRH6Z4Ug7Euw67Rf37IEJCdfXabZZQU7MmG
vYINgkCnapwb+niV/q5Yh6V8lZatkcC9vE18UYF1TwPlsC8A9oMDnkwd2Aax6Rq5TEaM3GqsO0th
CC6moz52/PRdLi0JtUab7a98zyNPzswYTXl1usv5eE9YcO0LMKAB9z8COo7OyIsW54Cb4pMbb6av
EICTx8JWEa25bQsiribBJfga9d08zQc2nGsWbnUo1gEZjFdyY86qXcIjTxGnlT0fYRReRxZ3AApL
AxCtY4AK+JkNDzBQMeYXMqXsWd/IPQBWsK+0JZ8cOhv61sM+0WFQa2JQkCaWm25MIFgJef02Dq8m
ANyLcR2kSnps9ymDyU7HRPWpiRy1eRgFRL30U+ub8+miM4Ul5XP84gElKzW0BROPTB2UALE/NyFd
bYErGNQYFgaXFUsJ+Bb3rIo+MjUUW+x+gNXpfya8JAtanklKWPokhzB1EeiCmrZADgy7dOCsU/qb
KJPO8NCJYvXxQyKeC/1IjRYqTlVDD3Kjqq26D+DyQFnlYuMJ7gZQsctKQeeAooSVOA07Qp4LuSMN
wLvxMx2G1F9AlBt0eGrrjHhv5+bTZI5J1MUnQMG9wf5OBc9lwnMSwWIm9aLZr+osrcYu9HjhbdKD
cyM0hvuTv9B/NgLrd4ksKFQhfdbtf8tbMEK9nxHqjphdjl9MJ6xYBbwuxUF+ezrWLlAJGFNleYHL
1MXl56d6WGGBLnB35cKuKf1yufgBPtIFBUyLNueZWaj7/Jr4j4XBE2sNOXsLigNvV0poUlmK6UTZ
5pNONAxvWCwubm9Giq4UMQyC9aP5fxEsyUZK27EQ2OMdHWjB26yoc9dPUKBZqvnWk3cGfPUOd6vW
XY3ZRo0Tzhl04CLzhP2oA32dKGImDD4sPTlkRj1bIasm2vtEXapfZCBnF9NeukeXsmk/W4DWu3Bl
Gdx7pP0eOvnGQjWsPEd91ZpaozBsoq4IwbS1H7MTYGR31NErhq5ribN5pN15GHU91m1QQjvv6D4y
WZX8UV5JMUWwLDDeJSLHXrVkT2CVH8/kIhan/kbb99N5lLjrGp8P3TNGVWwqtQpsk7TEgf2EHQW2
T/Gz/bm6GVGCBzbr/6Ssim4r2nbfERRpVgfjvtU+xmEGvXBSPoLpsGdiSwQN+LwEr92ymiDOY7Lm
pf2lSOZ6fL62pYxooCoAAjwl79DUbIoMwzCEaVHf/ZGAx7U3KVxpJKewqXKmn4Zd30+SMujSkjl/
WFyAuFTwsgdgceiucquYCzlxGgnPdb8LQzdui3B7OFfBUTGnWFJmjXwBbJd0F7IFHEHmZASQ7B8H
Gs51dPW8nkDjBVXK48h8Qiefr3HMZQXCKMyPiGafeDgHB0RXFvKqGss371NmMRWkdCtK8BgVSXHL
Sj1eXM4HRwFcR1IHCBfpkXdjkeZgbS2+y6+9GJ+CKbSnAr/RwS1BmpzFQWdZ1zt/uf7XJo3SlQPq
ZmVY1dS9SODEfRcdqojRAhsWTiLZlB+CWz/mz4+wlIrD9IILNeOVwQBKWYw7WiQZpYTnFIjcP7dX
Df7Cp2KbQJuph8vB+m87vlc/VJzx3DYmZHM1H9XoRHXikkYWVpsxtupH8xgDPgHQ8d6uPib82w7H
6ABiBsRa8rjPN5ewviVWisI8hEn2IwKsmfsHz2AK6RTQ6YieCZe/wO0oV+K1viKf5RyanlrpoLru
KAaaO+R+S6nCswVbIrFw0HHvCEZeg2IXqewIZgpCbBIzApcA/qRE5tp7dBxr6vvV2b8ezEodiXN3
lYtj13CE1iIypXgoSeSDSqDmH0Z/rh+53r2em29uYTKFhVd2W0wzqIYtejDG37eU57LAEV2/l0Cv
3u6PIGeRw+PUewoWN4T/lIm4DhaZe1Mxur2sBLzNOThcpFqHCF7IRCa5evpki36J/0+tRIU1t7bv
r78+Iun86YbMnNp0ebbd7r1ccCpvhngDC78fiLq32K5hnpdw4k6QuCJpantpmSsrWyNeL+bkFfJE
ajW8wZ122NO4LUC4gHI7oVErNkNhn2UX5mOtKwHyUB5Nrm08CRCdb60pFORph/S5IPjGTjwUv42x
LZEyE5INlrYvZqBUGdzUrpOGieitvh48l35yzAXqR+nunlV2FKHQM3WhRIlYGTzNDKguod+sDeUK
x/hSkg9Ir//8NXgqqVzR/4s9HS5OxnL49jhV3hUaYl1GLxSaBba0MCIXFrD+05AoI3g/WE8Vq2Br
PzZCVLOknL0IDs8vaLpUr4uqX5UV2F05vxObe4cHT/X1ro4UXSqwPYrbSMJHWsDg2odCVY2v//zm
yBVxVlNIhLRca7VbOAaNazMVWfivgljotPK18NfoVTEWFGzdPTbaHBDtSAcDsjV1BPIhpYkxH/Lw
vQVcO55eoXRMtedRvfsGo5WL5fnhGTtb8EbbfyBZUKiIhRt91NbOMfyPHgTJQl1CmvHgElHLiqdW
P8BBJRs9PWrhtz21muc+gQ2kuHyCGTg7NJHBvWBeHzrHpFpXlGoa5gFPLRFSztF0HIINUDjanSCd
Qj805AfMbQPqM/rik3OmfOkDSal3O2u1171/+hazuI6w5OVXTn9555oWolQKZ648MeMiyLZX3nqL
1njGIsO3ZYBrS98L9Nv3TxdVQZicROgrsZMwGlFx7CnX7s2H84GEKgUDRM94N6RQU4/KnkVndv+p
TSgP8Q5uvaNBwA0eLv8NSx7y6SQ+sTqlrEkSvOvRClmUOOEtOFzSnQwCYs9DYa8+IMr68vx7Wr49
KdNIKjRuIaxfv+KjdAfCrZtuiBM0Yty5SPD3DNUTQiOpLz2CjWJf3/QEA5qECV5xQrxMT+4uvL/0
Icvr2F7fA7R1jhT0fMRSU5UDqC4Pb3hUB7gztTfzLbIju0l2ZUG2hwhajbxuvv7ybiWGDrllxZz7
+p2gTMHvlwvuDs8CizvEhi3WuVY39alXCjaolOVNnL2jjTrrfIJmYIVfmOo+fcRTVJIGJqduHfEY
uzqruBRyQrrF2VTmlpBKESrLSMmob4ciaRHCK5NLeJOwT8i5QSW0OfGxG8sZhixerpoAVRVdcL1r
rFmX772arFM6/5YBMf+jtGmQbDBFERUnVmNR9FyMBxuaebcmB2jdKSbl5Os1+I9Qgr3+w/NmATv8
DMzJjXoPOaBV3CbCVWZ2Z7p9c3cYPUmLlMacReqrtxoZso4hb5i8KJgUM2IMFcbjFTetgkGG8umj
o8Jh6bZCcxuRqUqOSNj35FGzfOSUz9pcxyc1hr7J2wnN8U0sOx8nXtEedV2t7Lihy8M1YQBGTKDc
ZhEus6lF06UJtL+wu9432cORRbFNOL+w6NcbFrnXc4yRbkuoxYwkabs2Sbn5tc8y/tbEVZsWFBBd
ZbC62QUt48yyYW/BPTqtvDACNxkh7K/r61z8akAeli6mJD0Aacsik88xRv+4eVDCH90lIAcvErcw
UKBXrf/EGOGMR8GfHykeW4FBxAt8b34GKcqxgnbs4nKTVb8FgNzNp1S+xIqnr24TsFjDOU1LeGQn
nslc0Kr4vBCzUIUnJHJFQFzkIYJUjkYSIoxOgvcvDhjVsEVJTI6hXYg6Rgt+sGpG6lxFYUzz3cZU
qT05KL9R6x3nuf60A/N69RuUI7HgGCA0a5J05aefQWU8a49H3hpQZWd1iNGvFoSfHyxxtc4raTmD
/EF9f+04F5brVSj+FSLtswsSLYlVUsRU6GChy82r+0+pJb4LVFZl8BBLt6X+UNrUabsmQeMboMF1
7iMpMIgc1faLJmVII5EFjw3XksGEGRHQBo1GpTg4+0jVcXWjpus69MurWGVyA/IB9Y0t/r56oaxr
2MpW5URawMr5xjEYG3d09gY1h8vvC8//kxKyPbt/6mDaNjhR2/hDmjV+RIXPfXNMCiXgnvld5EAN
ZG8lCb+LAIlRasGoYVkHC1dPIhlElFcaEUbgQDrDe7a/+IEE1DDpS6GL5KdEuYFdA+UruONDCyCX
Yg7vibGhsYJb63pkfhQr69G92E4iRuAKUCmlZn2mi+/+E82JsayPazhyEn4q7qLEiPWuNrBDIZeO
49t6nu/SRUi9qr+w46Peupv4Jmc6mzCGSxR0cMF6g70/PCo4SrFp6zxwXE2TSE0swWgCieXglQiQ
COjmttOYtevJgRN8broRcBCp8Z5ty6P3DL5RNm5SqaqsknqrJ1qmAM/HtSl6Ck9BmA4Byb7Ouzy8
q0g50rNPDST/MV09vfWnWimniCoU4ui7G47K9McI8dkrFC3A0FX7ATDJGWqR/r+mhmkbKvozj+O5
bY9qO+YNkRAI7vCclTK2AU8JkA1Mfv3SmptE9yvqDHWZUUWHffTyKw+KypsumJjcfZb/NWpLIqU9
nzYx9ky1DltzZFMa+dFK6Ne2wwc/NvyIgFIkz8ln0pSeTQaJyTVtVyM9eRtjt+QeiB0lHf+IQj/i
7/dDMlCCOwjTp0+2mpohcBxEU0jtohnkDIaKl/hUvHg97AASKlDrKyfk5Xe0wRKAqgTBoLk9LFyl
NIGXlKvLs3lVzaTXcTl9KKSb/x8i7zU2uoctWh1VQMSPxTaLulvTD7/GXquj+qyCQ/kFp3ILyiA7
ssaovwmR3yczZb300r4n+nvClg+7VjMNwVuIp5Tee0kCqHRuMcj+9Xd1Mo7wK60z9IcZNEN2QHIt
/1qD1adzanBnirqpfzDIBvpgRs6zT+cIxXCYGQlkPSz6kdmCn8bGqdWz6UOdWST0JxyVjWj/Dh9S
70ESsh4cDEgpQFEcM0Ioz5oYd6ItJBBcwPxGK+YADGrDUP3M78XH4WZl3ss+GCn9+bM+dNx0fnA1
7xqSlhy7M4WmWMj5HPg8wU/pcYxMxRWrByjXW4cg3Gq5lduu/EA0OyPReBdjIDRECtDhayh/9v5J
OvXM85qnqeasFHz3HwZHj1nAHKrj5ZSyl2awPLh6Dx+ijUMvHjLW69yvXHLIUr3nETDL8bairHIZ
iFzwWn/0t/hw3X2j+mgO969F1ssjGRagQ5W9qXnuZbzrYQhNHpQkC6iXXHg7iWUTaNiZiHOjxtOB
VXWVX4Gv7tuKQ0CvvjznB+Z7Dj8qnrq2nVSSbSXyz8SwUtM+UgkuDtaR68NV4qky/zb8rvCZLtTE
hpTFI0ZfteWKjWFXUDZczGrgnmlbdH+NTG8iIf3oPdR24gwstGjADvDyEOrU7sYZE1Sj4Jekb7am
SrXA4wAH2A39AGFiGewDp1ggfaPH8DNb1nYUFER8hvAIz3+bdlA4ch+3nzxmTZx0+s9Cac3rbrrR
Xr5z4wivcQqSKjwicWcnPvX7QaVujC8QEhKj0Mp+y8IuZ0sRbUjdrFu6jQoHt5a/uvQAQ+HdDk6g
YdiS/hP1RA+7NWI0U/vfoBWhfHSuzGnSPlLUXP2iaS8L+EgZanU6pzKCseZdsJkrDuzSRaX+zCSm
l2LbPe+jwG2fcPWCJ716i1/XPlX9Unvs2Pd0fj2VzQ3zxlrlBtHCQVEF6nl+Rk49WuZAs+6winOR
WL0HvC+7yAgCh0iGfwMyym6l4+5rarr4CqH1QUx+Hl1co7BgfRBHhErhgl+j09yATo0B6K0AzfaI
kz4upLvzBwSknImOdjknydIN4cNtETGZDN0WU/RjC4Wtw7TqkvxqD9MFFyA1Y2vVFrPk+TIwpA52
0k/yWGn3CxY9bMS2mXuDAD6aSEu26w2ydOMcgSPFlTyBSxJT0UD2DrtVBCdPeOaqWT7hwgtKeNcA
VuuxyE50oCFSop2W9fxQJazI/IBaVgJ1JPD7AcAzWRiJqa4twXbGX2prBeStYfpBehL0pYQM3FAd
5kKP1VewGf5XxNo3fDTg1gg5A/SOCTF26XjIR1Mk405wISEghDiMrk+Cwi1Jr9nTtVx0UPA+C4Lz
0njDwrWEHXOAsB7Sdn+EA0TJar32QvlyxkTs+cJr+0fCaA8+nnyVjaCXQJMSTKHHCl6v+lo45TuA
m7qmRUPMpjGtLGP45ngCkvx/OBCWqNpqcMSyh63qRq5Phbp1aiu9Oixov2q3J8+/6OBbVPd1KbjO
Mj1Tg9VbIOb/zC2NBnuuOFyUoKSWFzkogAuLUi3iubzihnA2sGWK5lApHPWQ2Vj0gT4z3D+All/G
0UxLl2GKC6+hT0SWq8Qc/n/SIEeMuZ1JXhbFwaVmJNPB4gHJRwvbA6nQSYHmsCmVB8GETDG4bN8h
f0IAjRF+yukrSJ82eC/j64t6Z4GRDC7El1EctECPpJxORrfN9uvprGOcm5HLGJdfXUfDN+kvTWOW
aZkO0y8QX8X+v0LTruwwvqAXnaE+1EdeJyH7nIsLYO7vIN3E24O4mtiTBapIzP8eIfQsb+jaKdS9
T8ov6+sSzo9dtdPrWuSYoNQgotF30va1OkohLBgXJW1maRqcaPtB+pPvp0oKwtPpL26pG15L20AX
miojk5f7DIlHrcmta407saGDrsUeZcPHrG9U2WW9q3nHMvfGWTbqwunszB4Iq8hE1ULGMnYnr4gI
QEsEv0cMksr3hieqC2c3JAWd6AG5eYvEj7cVDF/gLV6fUfivu4juQncemeCVZWmx+1+q16O3mN/M
CMPSNIx15zeIa1B/xToDl0D2bYC/AnOLW+4u94441ixpc36HvVeOCYvdtRJYQCqLcrCHWSK3GQuE
xRi2T0AU3O9YkKtMEuCvR6GzqAMEPQF2ks/P+YYyadv+04gCPGkn9O1fmGgdofbbVTAlUkuuz/Gx
gd+Pb8Wp0t9fJqK/3/HH+JRdbJPDdPmBtGVrY2Tc6OrPP4MNCLy0F7gQdoWNtG+KLYp/kFgATzKB
qLygyRin60KztqsneSwkbi6PkSdp4p4zYdV25DV3a/24YUShwEB9fjnFXLW/agzv9l29GygB1OSr
12dhaXltSQMHjfRnVFm37QxWpKoKmPh5M/DZUfT9Hh3Y5OSfYk+ucc6Us3zh9yD3iJ3NAKrAIrEc
GsYljOBFaY5Z8FJeoeSyLo7yDTCfATRhzgGm5W1KtlsVJAyCcq5SJY3AERXTbkI4rG/baCRV98f4
fKqssYKdevwwVeWVm4/EEFugHdkDKzBqeuAFUpG+qjRTcTg4uoBqNitx+5HKFHnVzotuUMEBggcr
q8UMmE6/kKPRcEfwo3rXqHhyEwTB30aB/AEQWNazKeV269txo1YRgqjfKMoVUFSLq6ZeIQYF670y
hR5Qu+sLIUePWSKNRhIW0vhcd6HotYgS1w7dg5+qCEB8bDGP3nvZyBUyYuITZM/BJWdvUsK8QEDd
4ORbeAcXfY3dG2kbjBNG/NPNjbskY9ruXPrZDK/G//508w+Xrpv+5NDQFtCdDnWlPx+ig+wTnhaY
zMDw6DEgOTLvxUaVTU62sk518K8wE+dimF1Pbe1O/9b66HyqH0OPaCaZx/zHlN3h1uoGPoGlwekB
MoTZah+8fod8lwPGrlqEZZ6t3KiMgSkQLXuXoed0upTyDBWanndIOh4IDFI+l3snULXU0QnvMf+n
CBrl/ww2GlNbJLSZPMfIIPC6uLe4b0ZaQfFGzH9lBuifapCkus6Q/bObZnbVhtAapoArWIyjWgWQ
gOELB5qFaKUmzoddN/84nMS6LFlB9uRRSpmYcOBrGTlICrzIfDSJVc8dLuKjbekr69r7TL0fzdCL
aUWpBZ3HdGcRIQBdnTXz+mJ0Bid/irZzXpk1kJnSIb044pKN+8WJnhgk9Kxe/pKMlRYTXIQX01FF
+w1Bq0rjtFE4sbH2miVz64SPbAB6znl4Cjq0pJdIvA+Lkxox+BZSsur7o5KtTQzkJq4jdDXiONh8
f/0+5EratY81ZqyQltlNWAASw+mX1egHBw7p2DpwnMfawq1gIhtePKXSa3Ogqm4aS5ODAa1c0y2W
bpKL0s7uLlNKKd3HSvHujxL6KoBD56QScaA69ingx3bidwPYcUQiehOi7eLvaAvh0+da3tMqcvNW
JFxq85IXvjlSPGpihtJ0DsbGeAt24TPLv2uzWsr/w1yoVDcncNIzUN51wY4dzpDqte5Qe2UGMKqR
jX0IXWFQWHwu5H9U4wZ6P+MWAdO10gHuSijNOT6lN0HkFfQztXmBfs3L8jA2j0Zt4no4U7Hs26aY
FD1WUAY4JBojngPrHIwvH6icJMFCACqoD7/f5DF2Ys8SGfI4+FB4hoHwhGD47/cs/9oAS0In0uPf
X98xT/LF3Me0/Xt63YXJuDpSO4x+S2r6J2+lT0BhoyJJyRjRpeOCtjvjmy2jwcrtIH6AAfnb8V5Z
YEUybkt0U1yzK1WTG6OductYtVPJ+9rlx7zvmrcZj5l5NxsBMK3wCVFQm8SGPs9HQ2n6LKXoK/e9
IPc4iLeXsfsry0PXYaP2loZyA+s0LTTpcShG1fs4Y0Mi3qQXviyhagJeIPJ70m1YFszURwNtOQoz
swVkGd0FDSbO2/+sIZS0b5/AhZoiuzov5zASkeHSGM2lwrAHXVvkUQyZhkXFsILFneVq9AcchUgY
7B/XA0dHeCgNRKAlhuTYczTlSm7/4o2G/AILmCwR2bHkCjWa0V5/c1Yz6nNmKe8SQfIA0+WdEGyc
0q5fBBtoJx41Vir2QG9xpFgFHrXkQCEOIRLkwxavjY379sx+s8dxznNIYHSCWphT/PNpEKMf92Tw
3CVvDx4lVwwd7M80mgKgJx8ISVakdZA4hd0Iih10ZYNWEh2W1Ibd6exow1zffHRnbOvjPSQzJh7H
fEN+VClsqAxy1lIXSqrsBhs+iVGBf2/JkUMoQRMiFlXNxkSSkCNRmpB46m2j+f/XyTMwrv4YbX1S
o9MsUSZFYpaLmX6P0CeW7bN6spMe2tLaYuyGmq79TAS5wtvyZeWHS7/+XmHSoZyoWTsvjEECNfsQ
JE+wT8dInwgJWf1RduPn7fzaPXbFID9q69lO4a77hVU8G1UZtH/8BgS9QUq/qW8Y3ovvBvh2RyTN
VdY/lnyR7hLxNBHryFeCdequ0RFKKvk6AHOmwjM7mVRIyqbGDvlB6phuftRJ4uiHzy4sTEpq+ooy
zGSv3l6BenPMdrtBd4MaDNUoSQ7Ys/BGI/TkfGy5idSYx2Z5C6E6jilr11QTgySX9KHRSnl4uV51
hW+CWciVqUHm2hM4SLdEkLH+0aN066RAsS+ziWmrHeBZyWZWDiiE4XxJp0Wk0gEQesCtuNWq+ZM6
pCGOeGsFAzEeGfDnrItyGQF26xlx+c1EVG0ZzlcQi4HA+TYXq4sw/OeRSFZijzLCH53xpTciMCwg
5KNlkJOlgipzglvxruX/hWAxoNn/wBKaEsBpObpPaF1WsMsBnadBfyEo9p6y9G1kFSITUhTz76wz
lRRBoiR9e6H1ollwlobQZht9NWakDKTH+o5NMta9lBV+JcMCBruAK9JmwvlWj1FzLQn6mbEaBEKM
5wwqBI4+TJoVJ68w1E6uW2Nbl0m9o8AvUcpHUzwwd2KzRMRBVW231J8YHHlknJ17dgdvJqsxAQs3
QRWQwxuDQitfGyOskI/QkeI05fbX+kSFFIT4fYCSnUJaIr9RFiOtCdMWVxpBXPo0yT04hj0p07pk
Ohz+ZhjVCRGQtS+6MeaCwyr/Mb8pVCwHTMlh45xXselClXvhSQ5wJDr7Ua00T+cPYHFGt5WihfZc
ZBXPxf91cyhyrL0aJB9y7o5L9u2JAdbXyBpdEHgXHxldQn3ugCixe7AOu+fegUEW9Q4gX9C0nAPq
7zW6C0scb9uLzYG6n9cLTUmP5z+eiM0ruqC6B1WJv9bCK7u1BsfIO+Urps7HIHSc+lmM9YJcRX3d
wwlWQTO13CizC5ortSh6W7b/zMKjY0NJPTeopugNUuZyd2/l3yC2Q/S2TAOtyIOZEVR0CeCEr6dW
vEPpI1Wsta1LDWzbCYHgszSplJyy0V/4KgV7BhVXjKDS369ixywswpmMK9uzEPIWnMtsGq5VW3WT
BoYsNSvMUQqNcNHUEEVYvXyJuCb5tBKbWR3K8ePw6LDnGP1/dcps1k6OboOIx+S1S5RdhtNy+BwC
K2L8tTGOqm/qOrGkmSELXva6VAtF+qbEiYqmcn+TQyzswx2BkfTqrntxeuo7d+jKyo411cxygcoO
aWZRXc0vT0drgENnkzLH9fXY7DnVG3wslqDrfK6CYRYxK01xajmqi5kFQxLPqHYaAA5oM7qb9i6L
d5BeE8q3vyR4W+qSP7bECcCsWVPk0bud6+GCJCuTzvmVtP1UkEHFn4zBQZbCf8WkCqEWXzgaM5+3
KvurrlQmy6LfPleLHaBSaIU80aFTSAoyZo4eQ4yO5s/6+iYB17i0agZbcEnzT7kif+aSdvqTpW06
KLoIF7FLlYIhtGAZ85ZqwjJjiyZKzHTtAl3yrxnpczvBvn6SrIv/a3CVdTMtSbZUOPnQO52PskzB
qm5GgdKVuaeUzffO+WL45WV/xnsKGSsExLYbrIVHvQuhsF0v/uPndPaUjCwUTuRyK4ZtwiGiIFPT
YlT5B6wdyy6AStSPGJf58p5txt44cyXQiJ0o4HquL3vWLpLsUWAV1kKG0XxYC8ep5ObMtPOXo6s2
G+dunHMrx5I9j4Eg1ha/BozbhmM7Wv1AgtRKz4NGg9oAL1757Ln0lmxYkbLfQZLNZf+gV2CkrWZV
1vu4rFS0w0TV8At0EVCQYDCQUKIStlg54myxUQUZRJqRFUqeWBgPKx6Mu676VdDg1HNydNeUeZYa
Y5e+nRyJHx5fVVSJ3aOfDXR0U+I22wc85GkeQ3PhNW64lDQnks+FDRKeMuQVKudq1FgK8V2GWnln
r0Xty8uel1WBxbsn5cWuEYeNEcglO7K+J9ht2fgJOu9FF6IYXg+20THYLWuXIMIb+zP2e0F9QKvo
BBueHwgHMY/tANbJ/9BA47Vf4LYD0Or6rQYiIWoy0C4P48++4qIXErPgiAj9nsU7J5TmlALIFAEL
MybUTGE5fUcWb9p8WCyQGBNJ9OGPMvPC4FljQE0SP78Izc+5/mDSuIc7r4SEYwx7Df25QypogcoR
THYXVij9EyxmGXm5KZd1X2InkRs2Jb/oghvaii9wWDCrkYtsl0JXK8Fkk6ZThV/2JXVBS6twLo0Q
+367KNJP8KBcN290Svjc26lgH3lM1B/aTPUPazLhcB5QKp0EI3L7B9bvIUhUpAtI0chNgzVdPXdj
woCpLz0SUda+F8wPt/IFY7zyaek8waQAUszTQHj2CGJIEmL9BsrfZHwhOmZCQk6oZSlccYtYuaRa
ZhWHlceY/ECPRwUQsv6iEun3JTPeD46j1+RiBu+bJhsjxsN8Ky0RppDKl3bNQwMOSe6Y65NZh1Uh
HUR24ucF/rIDjOSfe+nL65f1gm9w1sGftKNgQ+tem7SKvomjet4XJaraUJu2Ga9PavjZq9RSFOnL
waPSPmzu7KHGOxyUGmMJxmqUdLE+b07BtnXbHxAohw9k7lc2ylEkWIivOPLSvbgaUCi8MV3wCDQ5
LnQCPGXIzbTS6Eg4OcGzqzhai54mtjnoNGWPqlKEU1739cKqBaB1sY8vsWTxcQgQ0lR26Qxt0GzX
E55a7RGVVV5l3B6G6FIoROjS0u3nfdOBeXhDv03J8QfOjPIdKUBIYQgswg2KFYDzFXNAWHor4Tse
Id/3Aq/TB0RXporavdUe3MSOCZG+2/TQnA3CNdzcc3CAnpWgBpnbwnXIMHY+hd3HaxGk8MvcAD1+
SaqwXR2GMfWWVuXA6WBkGN7N6YFw3umpfVTD7Ed+CouVv7noP8grh0f69IJiU6UIbHNO2TR16iNj
Cs9ndIsATAc/f7vvOF6VGFIAX93EnnpaD+jYZ+kRm/k/kAbosRG0OAzjnTdpRt1aAuQYLUYgULx/
6SCEiI+tJ4L922gDpKYzROh4Pi3c0Uitbd6b5dZbZI0BMmJlhW4Ex+JSZMP8CfUMZNu4Kpz/52tH
EHiuzZZtN1ADadmEgbdp0XH6PwgbeE+JwhweZe6kZ9spIZCebZFaZIIK7h4c64RRl4ORbpVy3IKm
lLyvBXHWq0VMLqVSPQ2d6fOt9iMjLs5uAYJJubcYO/vzKqQJHyqiI5A6XkHoqXT35NpftRnP6OLe
KROpDeJVk7Go5i3Nas4Vy7gFgjYzmyxo7s/bsgk6J+O5JS/CBuHLsemQM+Q1dd4P7ODz5xvVuGGq
zI2nXwj+QXUepG6My6TSz9JuLzXBBWnpEHWgwkCJeKmAS90NpQ2QcnSmpfIZeg9RyYZ6/sIaD8P+
i0TyiVDcWPZwggKI36dgQSVae3zqv8W9cD6urAb+hD+DHPsedUfs0GR4+iCxhVWDyPebZnvbDjsT
jb3UdQ74Lqz7Qv4zXh7JooL5DfbY37GTxp+L9xSsLZgQ0LVw3zpF3dx0AKcX3EVc4j340yfefJFd
R6AQNi3KvuGw924CXtPGSECbuZkwIKpwN1sGd2Q3ek3CtytQSY+RPbJa2PxL3RcsC6RYbRx+f9kJ
2ZCgaRYbQAeN41BoM2OhlPYblrjhSxhbfjUAns9tzss7Ip9TPKwQOoVHRiJ0Fwjawvzerg23BTCS
pqINPxLg30TzbjyKricSPaDvkdPAQagTl29OwKV5dyfAjV6oeq1F+QEkX5hQfbi4MUg+5GxpPZW5
w0GxrOwovYrN3+g1U58n/VjuHKeHj9aKECgi7SEhbKhJOG1tYAgWUMLxJpUw6H0tzCsY4n44WyVU
Q6z5wqbm+MGxRYEpbAp+Dm2wIDhKaEsZFxSuI7H9NGUw1cemAL6owi9oniKFs0ENupfFpHjAcNME
A4pHeE0QNmvw5B5dNayti0cjPYMmpm2p+4wCBXCnC1W0FgWGQU4U3iAhJGm9/3ghrv7h+iuPxhCB
vWugDtOwgnKM8regIcdTjRu9ZMymMSjEYvV35N0sTzsoGXBCpwJZPcUe/ByNhYI1lRRakVqOnstT
72C7jJtYYhGHYmastyrGTSemi5+A1wEB/BOXl2v0HFnJTVoFC61oPorf5CbsQLCK+BxyOpBNL1Hr
lkNdTd1FtRCP2MA9kx1tPzoNeHFJMRvRTkvE9lLGyxnQqMic6UvnI9BNWXkwIHI4BR1DKpwWMBmK
pVvoAdndrAckz29wyE3djl288cWTpp9ys9Q2Q/VSRRsXCjbW9WfvBkadv7gWABW1lCOYxS4FfvcL
QBAt37QRswu4WBVKjEIhnXCKXxXVoDjVxLpEiTnbPALn98NSg0tFWsPlazlaMtZS2ccFbV7R43fr
Iex3VWsvM1UgD1uXC4rnzwaFzesz+nZfvTkxGn4XkFlacXzUX4HMjNSII1NfpapEQGOkc7VbXP0S
txL7aA4kDlT9PS8Uq+Udrx5pSN+Eg5ddsur6Cq+mdej7JbqZiLQtl6RtJBBLtcNppcAqsAbEtBjG
pQm7xMdF8SXWweALEHjWmEkmn0Co7AGOUmBg0TJNK3Nx6ZWSHIKdpFXtzjB6dFL75gXbc7plvN0Z
6KlLgz9Wak/KuCifqMFinO2nivxYKhymmtLHp3hUGL3AoDVp4ggPK8mCXp5643xhSVI2joTj/1yB
POlUUdTPNmq0Ipn25RMm2LkqIx6LUaEUCGabHAMjv3Xm+Sy6WiuQVOKSLqOI0KKbxgH3L5NpITME
1MIA6jfaAbTkA1emB/beHZs8JaS3AT/QcTf7vmJQUf+37lO4hI5DQyDt6YjNkS+WVQKwPkl0uOan
xpcZ6dWn5DwMdIb2raGmVMupdjKxpIim/KNEraq1NE2WpbfRPLpcu6zrubB+E8VXJVMw3OVn9ddq
+d+zuXWCx7uwinBMYOrhSW+l86r+Oa64E0KFuYjqLyqiJMiYPF0ZDePXfejn7OBN8tsCpfHp7+Ba
lYCqGM+dAas6Emyu+yHQDPtSjGPWGF6puDPVeUrpbECndRn3I8L/F2dtr6dqXsIJhqyLck6pZ/zI
TULwLT6V6bDuJoJDOOWNGmI36GuYTXOY9VsJBCRxksLHAqKq0OlyEXT5iGRYPxd3sIhFWgXNBMnS
3PZmOz0G7Ko5br/pGKpyNMMy+YInzr0dpdqPqVc2V2kDDUvtASEjT5zjIKO/CE5u1zrgDRqh/cuq
ojxgNUe5zjbGdhSU39Hd84fjoUC4qgmJ7YxCM5qdNdkrjn9Q8cKA4b+Bfnzl9ydjguY2OdAX0cuF
PAeIQT5RLujaOrbHIL//i9klv42qZSi8BJBzbJImOuXigAen3eqsg7Cn9R/idAlyd1D6NxCXxcdT
MiZ0gy8Y9iC8cZpp6UfaafDmhtRRsxK0l/26Dsr9q74oXoXGxI0kCIbN1PH4/czmEwNhB0f/euuZ
rxZKmDAmjwXMG8JYffnivCEXSkqTydQGjUCbGvQ5xfRiEma0RcfVjcV6j3Wrvww7klhW8QcUbd+t
vpkV2GHrMDfRDmZ7nH7GzkuWZpCR+XUcR1awej8XWaYArQ0wJ971LP6h1mthvq3sXgqGmD+mrj9B
csaloPEX3PJNU9r65s0zkR0WQEGb022vOB2CoQCsRO8dvWH2jjkUc8nYxhXHWe9v+IxH9ZFrlX70
7dWB2srJzb3es2h/wMyP8EcEGMjaGldPZaZzHEb0HbTjz/AKlpGMHfj4G8eoPOjfgdcW22hsZYnn
K67KsIc3/2IpJY1mpMCuoN+s/PX+IhDvppLwZpFWiTAk/OVCLusStO1OJRAMc7GjcEubdqi1J7ka
Zba3Z5fVxClDZdRFi9dFcCp1NcGhERBPZDx4QaeFtjxBHVQ7GV2+XBojN8NJljPjHP/19u2Y3k/I
1uPKXIo+xC/+QWoPt3L7/7QgWprLxjgpBNkoA3Jw0wAGh4SDx+N+2aXi66uCxgjTXcmR6olhyNQB
5tvud6i4Q77G8WAYT8iO0ATO0iKGE5D2YnMwL1CT2uwbTq9cnYreyoJH9MWPSBhaz7lJbsnMm3fw
AbcrKFEfWBPUSxUA+98wHvqrTCdteHEqm4tkLFF6wB/haBLOuPRDLq5WQ/dOvtzfKLSVDqYejLxE
OjHEYyZPmgY35v1uxcZyJqy0iLQTS3sC8403axO7Yv7b0OL4WoYFerkq5S+Kl3XYEKJqnr1feR4l
F5/AZlinGDng0u00DtLi6sLT8ADuYqT9Ba5XJhKEUXSHPbC0auOMWc0DDvm3p6e/TEdclbOXjXXx
pEadqlg9/3/wa2t7/ZQKEWGwtGXh6cf4jx3NBwF10WU6oeiYRVDZZ29nZkhVAAxkKo/6+5nu9Znv
SwN6/gkj1NXpvkQvEf2zb03sfPmF+2lZMl1TXAzua/mjo9JGbyGzu9mgi//UlExl3lmxH6+bfsrm
T13VjPOCG24IVTaI23Og9PT7gFpEigDOdzRMV2D7GUA9FEJKHbAb3VXSWu1i+cQ887tYXMPq2e3A
3iCmVUlJ4iVBFxgNcLJXkcIC3I2lTIVqNOPGPH1c72o6z8CZF0sl9odTm4HVdfeMKTIR7R/Afo1/
7n9F5B2cFwLAsl/LqFoxOpwtF9guYlm0n/HgX720w3XKnnB6g/nDBUZYW0bPuNTjJv5wFe/4GoVu
FGdtycTvR2RwIh/LYWORfzwW+ANjBQRVvxs6nyzEol1i/ckYfn0yaqxLGI/zxXz/SXCs9FJUWvow
/NSGPqUr5bnoBOwbJxy6ivjtKIhP/T4FfrA80yZ3k+GuFWhjhDWRbWDN1LJ26/LMhTCtcl2savdg
Wefi0IgmHTv53o3xKmgatN9dolKy7OGsSFsyxbDRvY9kYGK1RydTVGzqTUUf8j4vMF58JO5A3VT4
5UleGJ2TFRgk+8KOu7E2Qp3w+FKGSUMUkhrQlp/f5gdVhZVNGcL1vJRhT/P1rrqUIajUrd75vO11
B/AnglDEuF3McVskLOJvCeDsIRA2DXpKVjOX/OatFIHKUxqz7+WvX/optGHpIzECIiQxsjp1OVV7
76L/51z0OizD08qYhj0PnQx7ORHmEth40v6IxG23k/9zDc1WcLkbdyJstFnUJ06bnB8J4PuCwqUM
dvrLFVlkg/vlc7JbyMqMBRR0FKrWVP+QbCarm8tH9LwIsWX3Rxv5/P9fK0erxFZWy2DZWtoqksRw
6sn+pJ0+gC4+tTmOz8BOgcAInSHSVR4UmJkYari72pYVZcavAj/kNsdXI8NCxDz9bJl6T+z+nG1h
FzkCUwoEQJs7M4TCq11YP7YvzDFclyWYZhcwm4YiCOOlLMGEsuUzr6t5/RcHcfXvzI0FsxkX5m3q
LZsKrQtwCgSAZq/+8HvmU6ueslPuMaDvROyZMDe8Xt8QHjFJYvNZbLuiIrT4dPGJ7BCfv94VPkGd
LFJlXYRLlXGxon4wcZjkA38oNvJpE5jd8YTONP72z/DIyDti4qmptN0iYJl6biIZh5PKmX2VUR/j
mEBXnnAiT0LPXzr9cMl1pkiWwBokde6HAI1HbBMA6XaTPcTj225wjW0Dmrd3O+7/y9WHyM5qdgG2
75DbJwTDfAw9HQgiJACEumR4o1GWPqwttLBlJ/eqPu73QCoQgT2lxfo9wHTY7au+RkMJDzzGf1OC
psHwFCb9DWRpNl42i5juBST32ye133jo6hdSXzvF37kWTio0n9y23foYetyD6R0NB/1sMPvTR91+
toeZ+i7ppjKh8K8vnFETmqKRHXVkxd39z4DJujk+O5TomEH6YAa3Dla7vVtngz/dogYZ74Vtg4nZ
bo/+80JlMQf9LG+GQwPMvxOFeOy9MVrx6DmXhQYs5Y20ZF7K6DWQikZmckY2H/4ms7cjJpTSZZB7
6oXLJvS4Y2xDOSKlAflnUtBuTbJizWm30T5GwjbtvZxkqFZ/XLE/6wTCgppAlkgC2UPIIdaWQGM4
2Lqly6iuxVTbncKS91sCmNUpavJAXboLZTksWOTkV+rjkce9CdkTHPrPDzO2ZZN0t5o1tqA86DW+
vLidgkNK0YhcEFIBY/yCLSsbacOmBPf37cJEQr9P/thkYwy5NGSbI2P9qDVE9q9AujFpZnDsO4Yz
RJfILPYB2S+HuiZh1Za1GHsnZ2oHa5WpTBzcWLVqgfry3+V0BDEbdVY1nncSEKAWWJADTqfekgPt
DjT6NO6l4QVQU+ooPzz6/dlDJghI6ZQPrlliKWsjDrLZP0pyIfKyIK+p5iHdAxPSpdYrW0KxBuPZ
byr3yuUaELI8syVE723xTBUXzWjEspt+o+IcCrHBUfutjPrkAohXDUy+7bwv0e5ARBsz0d/3g1SA
h4k+kb0khnbJGgXcdDmPuUXgO4ii/rzIFfHFaaSwV3e9TcLxVWuoK8Z4ipuS7wQRWk+aoSF8D/mA
IiS1RtteE2btLd7DVrRoQwVNlZW96L+LLTimizpV3w4PGh12VIrpe2XhoVttKkIdBvoEGQMETcbe
rkA0HY+NA/GxY37ZujHf9VOJyQUzolkv5gEmTgR5wc0eXMnCjzU4sarlCi2i8Pw/I2JxlIR9EFKc
FMUaJ4RRcP7l0GDo3LQTdwRcuK+Kam7XnseOQajeBqMRnsvGhtT7mm2vXLxfnQyI8z+MvTPzEiEx
SGqr+66ZxBF/Gn5IjFelDvgef6fqMxShBuzwNim2kCRK4iKIX63U8VGqA1rUrI/AkU1kN5aSWG3/
2GEnLWeOCGxALbCZdVVi/7BXGWFRbYgoYryeHe42phmGKEAFErh8gGE8wV0m1szy3ZmkGL7dRBJB
gkf/1MSG4Z29SqGUbwLI+LjI/bHAiM1x13nbo63y2t4j+hc2nEOGL4bHHe3dP+qNXd9zGPJDjgqD
j2jWPIVN3pNrrpLQZ8Y2PM2SMkMXuMH42t7XveJ7NJADZHv0GAW9BmjJZzYaPhYXc5i+A/tR9G1h
lcX52QeVXb8EmJHI4pCy3QJ+aM7T9qnxCA2oCC6e41At308N5Hemn8cDCnFOxb6+VNg5T2mOWWEs
RDM9C/323Jr8lsZunwdBz1YruBObBDkydVAHWXd69HlAvl5l3kS7y/NoLzUPXSN0KMCHioNraLak
dwf+EAn6VshY7M5FNhUyy28E26iUJBW0nULHw1gcS58E7JZYhX7ej3dHMh8oMesRyJeqoCqEIPbr
fnu/eoe3gncu4TDlrGdZfF3v3AXjNP1u24vDWKcx5iB6ul/h4jrv/o5k/eMn+avBASZPF9a0G5J/
d3GKX3LetS9tcmVpgtBdNL3wPerfxIEL8xLRY+cj5IWBUPiE0BCpKISnsJ92ir7Epkf/2RWDMxsQ
9r0BHULD5AT/pPenOkRYLKcuiktXPndhsFggKcxt/p8VtCUD1cmx1pQaiQj6oElBdTlQISLP6n/l
7yZv89g6rt9fFV/oNTAu+g/NBp/HsNkOzMJ9ep79CibZfbXRBXo3AKC122swW1IjfdxTDStKrcC0
zaBeA13EmfNJZLcTZApcxSQOArJfgGbW1soYPLNkKNtr+L/a9PbG4WiwpioQjyN741A1xtVgdbRL
fwC6Y0CDo0+L5d0cecmcJH6qE0zkyPAR0Ie7JUnsMzg8e18wLM5zT9M0V7pAHFC4JFMCS5L5Ed8e
2dM/2a5UAKQKjUOctn9fbbbwsaFaV3Yx0WDyEHvZSn/LFn3V0UiLGJUJUuw3U+2lYuED1I3Yjxng
zJYvrk1AIDfvTi4ntap/B2yXi0mNkRphtT1B281b7icl7NxWw0TApeA7tqtWFL5jTmPlW7DLaGQb
DhFhDvBFWHf1Hx4iuvWcb2+A4tLaLgnWGfvnTFIKv6RYuhjJIYM3PHI2NiBOD6SAWtnfr4cNtvJH
bpR+g6n4fYfdt86DHecCCIFjBDNEIamfL/09HqRHpZydnJsz3hkFMhtt5Lox1LazXsCErejBHXWP
wy5p0uyJ1zVwKQLD8qlrQB2lSsVfPIO+qu4AO3Jaz4aVWgMhkAuecGzw4AjRy+2YVREYRK5tDRLf
K6N9yIZBJkl9YT4b5cEBjVNzvHHdSAuGPkmdqmOBTfnIDhQzFEeHjsBifSCAM9cRcn+DJ24YEdlB
ffMlE+EAFgCp+PXoTJWHKE3PVU8ve+WV13cIMs1VXnmjviuz8FBjUxnJsPFqHJGEda1ODsAF8x8u
p58ccXe3bk8OQxHfQwyMIab2KQ/5iFNs8jG+64fiLmXChpUj8Z9uR0qIAw2qdB2EP1ecNnQ1QXdh
RBuHxLy4bFcgWMAHU9QSffE24o9c+Yc8MKUrUmrCcZ6jZUWtA+S5afhiPU+slaz95OdgkdRZh37X
UPr4ArVtTyjgQsQ4yG4jvVsxQ4t/U4V5m/i/InSoodH1U7PVMcboJFQIjn/H/j6i4zlFR8FOU1tN
XkH7BlZ1spGstPpltXmJQDa7wDaO5gzuxHmvLGdmCrm0UNqD1g6xcfBkJipIvmrLTuY1qbepL9KN
+ewlv5WQG2fl0U2uTGyfsZXk5YW4x2r6qrj4mcee8kBg3qObAJ2edEnXNlaq/WWBhUeBeKDN+32/
1RNoumOFd0YocnTl6xqAlsSbvUMMrGpOD8mzCnDvOzIHA07jgQwzdPyb+dgQOjSc9q3QxHgSnd9z
IDM0LwOYwGI6CNFBmlpTK1pImuo+xyoFIJuyLMlwa6FlNv3hmWb6T+xUQjjNWU5Cju/4iyhjsbl6
8JpQKC5OWpUQLVF2RQUtteeVZL2h8BHAyabanQuaZr0xv6V98et26jip3BLUr2W/9tXbvj6FbPp2
25EinVD/t26+SqacEts8L21QogLRDHVjen2niQ7omfRGwVWsUgrqHSMXeMYuuzQDC3Q4S+H0eHZt
hno5v9Kf/OQWR7TbxbKsUWonYO/1oQWEG4sI4BjzACvx7EHxsU4uvQCF8xuIlIeRF7JEzJe2RawM
0JqkAl5kIaa9OPLGeMtdR89VxKGhRKCfs8AiKN5/sYI+NsSw3IDRc37jxeeiCZ6OLXGfjRc50Pm7
7O9+06Xq6kaE2UXpM2YiUgu3b/Ec4fwgrDlrcugCjlvA0kLi9hBgKddimoe7TaEfjnJBfes6gBAZ
AzwkgsjoflEqNeK43eCufz4afmu+CIVgdVXnrDqsukHgiSJ9tPlWpJTfa72JqRxEfiy7C2jRcrb+
zTM2xNMvCIAdZlUTzcwmM+3XQXiCa8Lws05BMo60pEsVYEcOh8ajF6jblaRUTS56hNtbLuaFbMgy
KOiv72dqZTqgIqz5ncGlP+6qJ0yfG9iMm/w8kiXLpBByo9QcYYXIHjhoTWXKmjNkOqfKYAeEs4TD
mebsq6iiOreCfvRcK+P2y1dGvW+H3xcc+Zah/u2jSF9XgRlTdr5/hTm4gGm0tBv9O/2e7YdLT9Gq
N57DOazKM4zKa8/y4S/Wemp/uNJWpCgKM1tTFroXo+9ccUt0LpSxFW0hMWbYkguD6cMBc30bzQo8
aDZWA/m3iG4bTms9cuy5NYqjshwO4WcoD5XzK4JzjqyOIUOEMtWaMJUKQBLFxidgUfVS2LFCMeZQ
u7mkrNDw14WeSEq/QAOwy41eKMW1PLSEIRvvhTXsiScyPAYS5zq3YizZmWMcq/5H3V2TgG7TQTlv
MBQ46fdNT+sZ513f2A7l+eZ735+hBsKiJSe9Qkzh9RqJlLxNBoUPfIOYP8obN4UD0AaMH5niN2V3
kcGeIbZ/x/+uRDRCmMPRMEUuKPJxWCI7V53rVAuSmhmYwrtobrsq9x6A1loy9XzIKI7sPLHTojh3
vHEvr8cISSg5n/I0n+Wcrv8Wvma/irs6lg8K1X2ilg9SUf9BrF4IH+cOtQHMGCSA73RA3KRY2KNU
KE+A77NpRRbvzuNEZ00b4keMn1YUsxR9I8dEQRcd9AudAaFWzCPiDELWIkMCjIv481ryHDUbt9yQ
l30TdW2eABtrHc4KJmzCf33xO7bLu5C+bOCPpSyd4xmtVzft5fX0x5yDvVTxGvqebfuZJHBjMEZf
z05Xg4gIrTtkK/AVgwnvLPNO8yM9wzfX+bjms6pJXsaU1kIan6d+FQclUtSsYRcsYvFNQEkgeB5O
sFqnSiId5FYMeVY6qpC2USz64w6fdTUNkAmTrNujlsez7BrfX8gSs+2pBTB4yOBgXzMLUN6DhM8I
2JtSrV5CrMnBfujPUsI2BuyacoV+oSeO9aPLDGDDDMxyud0iE2tMe7KU5sD+GtnSBvtcdyGqbOtI
pCbYkssCdU5zMnaWVMSDklUvW5usu1smINKYQ5rREIEKHEwt/bwvvef2Gh4r+uTTkjdFkDmXPOhO
3lVG2TDOgLp6hquVylpAqKj7IPJUMXoB0WAW6pFpATKYJP+54AcTIyUZM2LsVSMawdHCWq7P5ulu
xPqrEk+OeMoWrhalotxXnc6ARefuVJsvfnSktcLowrbF7x49PidxV8cXdsImR7gVKC2HKkeE+xFy
zkcjO80Lr9SuNP+uIauHLYkZ3z5snLU39GsMd2ebHAJm6ABLpatceyRVGGui2SN7LDzpjGjcA/UZ
LFlssb4N+y9DcUul13zhQqtv41GIa1UsFiTc+MOUOrJlHryY0i2SiHUSV9kJ4nqmaayw8PSYcW01
SzcrAY0JbhU9Wgnl+CC/KGOKijuyL2llUjiltd/VBUdnPFP3WoC0Nhc4Rr15han3SYzoAvTtEHa2
DsV550YS8NpC3lCPg0BXzacXdds6DT8x658Lr3pCgKpD+Pewf9ZAohy6VMyGI/skefk1ivhN1AHc
1lfw///ILKB7BgegqRhhS1sctDHzbdFDERyRzM4HGTRHdkkf1ayoxsxJNUvhr4jPk6keZislNb5O
CkRBNO6meNCqmalxDyYh9+cDDMxRxvPMK8gLyFPTB7pLLoqtkkY4cFAEk5u5LfVKEjFoR3Rv7jJT
SuXoDUIrin9HdKnpnbIwn8Zy6Qn0HZQ4AiGVuXdWfkVLIUjSSYAigyySs95QvSHH2G7CySFl5ZH5
xhRSpPQsqnvUTadAjRLN708vw6DBKjkfelqajIkvXLDcgXFR6+U/EdH0RAoWwTuM2nX5DSIFXxbc
O9JQJAwdT/9Jh7GGPytr1ZOFIWuLbAG8PMp0iQT4vZ/1IoP6CcvMEU5hF/Of4H/t+0TJvvkqCTtS
B/aEIx4HKDUGX23KnLemp72wL4+aHnxAXS6Kb9wz5GiGmk0eqqGumr8bQkgmqVbuiI1zYVdrv2Kj
xsogPAe/ZB6hrGTmebHUbrfq4EiAgQSq/rurdlv3h7K1VXFWVtjdTKo9wczjixZuPG//4VHKcdfW
nJty2Of3DXG7+HKZZOi64phveq7/YmFpTKKC7Zhv8941wrsgc6Fe3vZ228wEZjPWMiCyuiASmGwF
UzVUE2H8KmaJ5W/xkxg+97xNODwka/6S5HUxrZcVg7yBvIhhKs9b/ZlD4BOaKwUymUldVu5K4ywf
6omyeoHNwbr5rpuGNMUsz1Bjza+LJKrzZLNScSBK3rU2sQAelFSshRTvZHQyrRXQFXN3V6xZDO9Q
o+VOQB2AW7HnnAyDrCYQ3ivwkjmAF2bZfMJqnXKhKY7PQoVZk81mRiWmFO0U01uVkrF7FKJEXwsi
dzEVVjqcqIeph6G1QtoLM6aQHopSL0oSRJZoBVMqgzBNoKLRe5tQ5JiIlml8whWxMHDgg5Q1OEan
SjCo2Xu32kb85caXZbewoiojkPD4/Xvvc2PtkQtjFZFF2/0X98LChCFkS/nbT5vV6f1TxXCfmHuJ
49WidbVJf2Udck+808dLvc/KmrexNLP3swWy8quR3NgRQ5lTATwMLKI9BrgW1E17lIecSFyxMskl
qjRRD3X1pCGxdTvgDXtyD32C2q7AnCjExL5czStbU2rOqk/JPM8Vc4IJlljajVPGPy8o2Y45/iIv
PRkYlHpcm5s8hE4Bgd1hcq/yNxjDLjpCzaxplIQwwpGGlng4VN8evOwFnkGn3u1DrgHZf9EM8ZUm
iv8XUaqel5bdmvmS2XEMIWsMQJSNYGilWOFEm72C6PWpOrNSUgc5NEd8Rnv80iChjkM9OOUhLVo8
F+9PHJ3695heib/FalwYTY7ZbXGep/N1Y+hWt8agu89Zq3dkusjwDBR4Jc+sw8FgXAkqdfh1BcNR
rxJBw+bYa0MmxRQAmDr9wdWIgKNYwwqPaK/JrcdCNTHUQ88pe3DS7MZuaAcEvG66LKgbXaJSNnvK
bfPyQrl2yFtzOAjwvdoGVcFhFnyqkXX/t4NW24FSJUn6dzBSDP8W5mC45DC4oQYY39LOTGet1kY9
8ugC5G+wNku3HT4boutNOmWde8cripdoKSXkr8p1ZWrZjAZKtDWHavZ+XZZaQAhnOoXcSzJt+Pdw
QVIbeuEkepNy+hddFTz+2+5P0Tlrfk3+jgD4TZcZLQtilkQGd4ZQ8CPS+QG2XCtKI38wh2zx7sEy
+iCco/a7vU//CI7/NLRhH6exNbFGGzDH5g07/iYg09v9grk7a/ZmxDy2L5MtqBCVa8xvgdVz/DVO
FLx88WQKbiTZzIVOefoXOQmwdwA2smxb061NeCQJRHeK58uAxJejktg0mPB5CrH8WaV3VSuHIEhn
w3a/ZlOQ/fIERaT+PKOvRbMh9moVNDR52aF7DPNH8EB8ekI8zh6Vbl79kXfDOWCBcW+v8TdzU0qQ
kfiajFGLIus/p6yYDdQ78XXlMVUnBEMlaDB5Wk8Sf5Xx2RsWa9bzy9enUTJsinD7ZGZk8CXZ/PCf
zWDM+7Btq+UqCxPPQEOZmAraNPpBvpl27xHQEfkiAXv24ww+rF7o5GoDT4jXi3EPuyNPaTAniJat
u9spZ0NjIFsWbfg0X5sBUtlKpUimwW43TH/FQ62HT+Qv1RLCVBfi9V4XYXSBH5ytyYFOb6TtjEQ4
mkWJdBSSYjQEfSOeNLtTVF05jUpqsZ62ycC4zO/D+/dQwyNnAE9rRKKK3fvAlnK+TRimWBY/4M0a
J+dXk3hrWghUb17nwhYIKWKQDgCiEKT/yHYZ1TuRr6bERP58zSJlpTZl7dEvgf2WbT2WCL8EIhVA
5WYgte1QdVF1ILDR2Lqu/whuYTNArn9sgkreYS6TOx4xNbu/HpTp6zRvljXRLPgN2Ut41sud0vhW
tB1Q3PCPsmmzuK4Ua0azhkgHG1B9l9QQqhn2bviBMtJAH20yxSIjGyB9Tz36bRN6wDV/Z9MOmcI/
sTsrpjMsL0O3kfAP4zn8TSab617DEFedec7XDwFkiTbwsFLWrkL8Ww0+EyjBla15f4IW+Zr7RV6O
QFvKH1a9FYkRoTLJ0DWCyT25+YIWP1inmLBSDe+wFwjbUqBsTGwZkyZtZqRvu6HYPLrQpVlulM3K
PE8BwPN/ihop4lZOyS1Cm9yxWF/tvGHQjfPwTttDZM0xi9myrWHj8OVcfSkWKq2v+7h9f4HyNCXK
wj8YnD48HOHeSvfepAro690zCMT7f3c75tWXvArxpBuTrU7kgCUOU7nhyS83mFW9GX71EUsM7B5e
4luwTQRLDNY6BpItkTQkEwBn944nesoCkJSl07Bg5iUe3nZKXogB3gbest0kmARhx2Rrb4Kv2W5e
DyE8vzlRIP5ubhslL1b/q4mL59Y/nC13q3gDAuY319AbIpVc2fJjqaFowFhdME5LTYrKz0JeIEMc
gFLsuTA09Qo9gES6p+OfcuirNt7EhYZXOG7nP6XRsTDsAktV3j5coV+PeYi2OP1WOIcXWSM5iBlB
cmhBkhsYI7K8GEX7qSyLdxQeIx4eS0zvHjpi9Ybn5MLVAkK9HawgirGyJ5bKFfzsWgVDQYcngLbb
aq0MUyzJRAJ3PkGQbOmFFbseT//DBiRrhpULuxnZsq4v7KPSfu8f87r1rinwiB2/5ZgBgeQWKpp0
dwGEiQNmEErDe3G3Nc7tXgKQhRF04j0iDJxIWUsyWwkuIOIyevR9z9xHmUNaXPNsbWqfU53Awt83
1wSGDcA8uGKoYWTxPohD/+iS1T2FOnLfaxfDOynHOpb6w3wYpukVdfYoAQJuqg9DzR4z892Zplp+
GEhmFENKJAC7AIgXZNi1IuyjLBrmYIcTSr1TBSKMd7r4TOe5cp53ejlwVcU+hUyvM5WWPuLQlMTD
u1xyotBKOAS9AN74egFHRgTij6SGkP1B8CjxrdonTLEXiY8bv0mwLde0H06iWU7BBBtLIs/6kNBS
JplW9R7oFqn6XlrI6/XAbo+siUysuCAaDzubja+pLkYv7KPvCR1HwF/Q+xq77khH3h/gAHB01Ptp
Y3TrQbTIAyj9FTipqNnIv9C3uQchV5oP/XHsqbm8fbu6drCCflFNoSRshoFnp1xGWneDscSJchP6
DJ+L8bUlgTmjtPTm6408RY2OseBr+WhNSwO8bm0GnGVzwYPZrZg0Ctycgd+NM5Y0H6Jc3kwAXuxi
Svo0Volec1ETBOfZj/7QlFMUep9q+Jy/p2WXjSkR2YOPgdhGitM+FGlR38iRzECS+XMAFJixamaB
Meqe5+DBJRSbsR8p8iuRKC3qkKynEuC7kkRnzAycon8oiOfZ9OLn/JhB822nlej+OohQ67rVXELE
CdgdANdhmdJz6nBgEoT5tnPsyc7b7MrlohsFvZOaC9X07fmtm9YqK3YcTAc/xwSqsPDBUo3SjBX5
FRYVdJBjkx0oAe5eFLM4VVRZsVbvVyHYJHsF7Vh1Jlt6BflZSDGeTUBarqSJoEXCf+3Pq9lx/MWD
0kRh6wnwKx6Lm9c7HStzR+GgApS1piXrY6XPUFnkEt5TxUoVPw6qn12YdylRjNKyDNTZCzVuUN1D
7bQVSshZoPG/ysGGQKerbXjctpek7Cf1Rwlyq+jNY93f+/PLuq1B94Y3uq7VvOV5d98CGCE4PQ4f
xcibTq8N3UNI6//ZyoIxB6R9mQQdMmQebeefbn0aXwxWNSDbdVwBa+9QRNtqr5bS6k87DM4DFdqC
lDv/2c8nHH8fmGYyQLTs5cecIzHcoL9SRBqceBvgwrej6F0ZqOy3YN5pk4fmE6uysxdtwSXW8y7O
9lImst1VG2d9fvqqFZ1Iv496gYVQhcOM2fFjqmGzEZCm7PT2LOshXKsyn2mIRxDgG3ADmPHO7zcb
GAWsb9n5LWZhUe4BkhOfKQLzHYD8XUsZvhk6sg0lKJ7L4TSnf7Y7oSemXgZhqER9Hxa0NAfxUIDt
0W6PPw3MO+mKRV2QZMWefHDkHMLIXaIfFEk2mNQioimmaHToLAxEozdaRkTdyfy2yqTPQdtH2JPF
O+Dn0A5DpkKI+YGTWlyZCfuqlovZii++li/LremEf7YH31FXjxtNou8bkLS5f2dkmg8GCnyGhVtJ
tWxeja3J62BmxF3f1lWqGx89NodyFAUemsQbn0XgXGZbYa6r57yA4TFx/QSbOXE2FzAzu6vVlxPu
powd4vn3BYzGgEArRYu02KPvq/EAfP7SMPejnu6rlRkKcTT4NHAilYTuTOSc1okkhf22mVqJw2lH
ztE7O1oD1/D+6IPj1H0RBjysWD7hQDUj9suLxmG7S99kK9W8MyIp1tnXgqu+FekNYAyvXn22J4PB
7JPYjrVrcTAQ2dxWtBCU9kI1NCIA2mVtnYZ+TF+FdBD2YT27brWWg9LZZat1bDJNTiqBTPVzy2GF
HqGqb1dMR3tLGVW9vSIGLUzdI/zksbgUr1k0VFZeKcTGDBBX1o8hViLNvcFxVTFqBKEA0JTUeZ2p
mI8QeA1Is9Y80aJzijSOipoS4ogYK80x1xspRyUFMcJJ+4x5Zsnm8DpmcqwNF3VrXQjDGWxcO75d
M5D+a99VXef1+8+iXxa91aU0+aWT7i0Y/+emDhxe4zMBrApwvtzlKesvLUzRWzXnBU6L2NF6wM00
a6cadKb32ZenrU9UwERS28kOUKk84AZJ2hZ+2S+h2j4Gaaz4TeCw3loXwbFkmXjzg6Aql9RK20L0
xnhvbB6SlfDNNvRxzcT66hzqOt5fm1b/w8kw5FxEDiCJf1EnJnd+PDmX1nJkshIc38UhcSQAoFcM
BnRbg56S2qNNiaPuAE+IE/aBmVxUs7DKSYwFkn8cGtU9x8y3k/uevWLZzMpzZqEs4IlNL4k/lVSQ
pMuYqPYVz3ISUup50+c5VnXjIeDv0GhUbwPOdU6BQvW1aEJ+Jf7g+GzsTnUOyMVRjjT1kTbDHwxp
OcgregDnw0XZTwPCwWnrYp/kDoHfyLgVAtZo5Zjj3aijWJX5VIxiB2jYkKzyBfWyoKqk6unnqymQ
4z6vdCS/w23BH4wEjnudf+a9fOeg91AKIzhBujQncZS5QOstNZs1PSnQTOB9JRGFTXlSWwen5JwL
iiOTVtuP+KpWgSEyll6K2k2h5Az0gExztKfxFtcCawmvVFTZBHwMLKFEvcY2eiibSp9mJ27Iprn4
GZYjBa3HFp3TxYSwuWcuOtDeosHnE8iILXvJaSdkPzZB9CUIk/4tM4LsmUCh4rfhW1S3hnbERS68
CIoLM7RT9nATWUGly/tqSryvfHY0o37qhTktMSS9S5N2hP5ykHJQ1GCPLiJW6lCsqLcf6LgChKRX
OtYhTcs3crVbG/AcZOz/Sko/d5HWYqEXypyhvGLatDXqOUwGuOETlhnEUEPH8sPEPqbR3dXWIAOc
xm7V8kJZDrergvsQR8PEf6GZCi9uTTCavff9/IKeBTKkODOBbkBs0KX1hUHNNu2CGHxIZ+DedRmk
+ZmNdaKXzT/x/5GvTxZu6BXdWytg/7OfpbPPwsyVbbUkWupoGHyocxkjcwCsa9TRrJDam+Hfrs0u
vN6LfqzHXtLX0c5sSfYK/iSjWwDfCZZlTuDt90Twm+uSaz0R2cFLk0VD9tOWbRvqgcCIuH6PeboA
FkhFWG0n86dcwG+5vdLkr1KG3g4I7Jv+oUPNEVa21e7lBhOwVOS+TWSO6+r+HWyWiYq/x2Aj5aj8
gpDm0k8HnUIA3FNzUsPTbVWML3SHr5pI06+M8cHaF2jpwiSvzSz6wQO1iEVya9lER3bsSbXKMKKS
J+g1TKrTW6ZCqzjteIjfnQDVrsowISF0z+zcIkS2t61gjrhPKszVNs5GhSCEbYIoh8WpgC7c9f85
oJvjS+8X5tPJDD2DcqZP8cVjvbSDtQJZ/BdApBBCAnThGyrA2PMAxKEgXdGAGWkP1gAizawZS4NV
mFofYDBST5nh6HWy6kzJxy9w+Gpp1C0nBi2Sbik0nnxQVP4F8Q1Q4/i7iFd87xoRfgnRjQdRqo7X
K9qjES8/Lf4ytj+XA8lrkSqtx1qhXIFnY0zz+klCv6ery+RjPyK0g2dGPp8JoN7BVb6HZdYduwG7
k9J94DxSXh1PdJ2SlFRbe9DS3oa5ditmvA+tr2GIF1yiRUZ5ufSpJ2tdFPkRlBEgpXd8vGW+lzu+
Jr6sCogKtBA/MsPcmMZg6uwz89U1rQowPyQ6t+K/XZzxOAVgXJm9oakGhyF9wlKF2O/DSmHePWxZ
iIrN1R2NBDbPFc7+cMtD5oy42kOeDrJmY72pgVoTiNMJw8KKz2jzpv6QWLo9zr9Eo79/rlFHENiO
JLOQimBma1f269UqjnbNOIDP3CrA87GDrgD99ooUWn6oXk9AcqkcmhkPfWuzr7hvPPM1i6lYknFQ
+gVWDbhVbExHh3A6dVKocPUZ3rokhj09gdc8Q1mF6zoznS3wtYhyka2AD9ckJVMulbpaS51H+F5+
59bKeQOzUPmEVC82/KG9h94MoLnn8q1aa7msvI9KlXpDNfnOx8ti5LdWcFKmXg7FqMMjdTOEut/m
nhl03MKmHiXQioB669P6RHdKz5Z5mWmVyFWyLfEX+MTT/2CvLSbw9Zly3oyKfr7292NqwHNW9KTB
In2XRm2IKpXO7Eb4V4HJxrWNn1PW/8Amz+uybOCoQYYRuOyZMPmPtMFAO4WCAIMFM78l30a8zye/
KTE4Lw/nXljaO5+JD2JSY7NVmB40OA3VDVJHGxxR4IAGeSybD2CZxDpTW7AV155sCD7DVmWpTtWA
DSbm6oU43oXtN7EN8nh7xhj4LmBkWazTr0JvAgQ/W9DkQqdCfuwLS39vHoLu6RTZQcEZxJq40cxS
GxqXdlDmJtxCAIb4tDqdk7uhQv1qmqYkRAJChNca9SspQQbBG5AQ7MaVwBO7/es/wqcNQwbyeNNF
CuEAnzIwHhxCXONE0GzNvmMQ61sIWA0xvRGsjx31oKTVs4qmrGYV5M1sDl8p3XETbWdZMjrxuxcD
NeLX6jmnalAREi92XNvoZ7zYdPWfN9kRjDivQw+BwRINjdzN28pKZTdWd7upi4llYGvuu+fFrtQw
fe/0CsDTjOg/M1VgrVfZ/ODF9fqElsqrhKdojHSUm8EPdcKEClSbw+A/WYQqgl3vjxU2gkBDxoyq
ZiM61JuTnLcN1AVGVNgcjvNbqS6SMGvwYkl8EkGhEwT7xbqNeBXPP0iXB1VH4GlNEuIpT+9mwV9Z
yj8vnGlJPuYS34IkR2uOhINblkeRp4VXt+rp+IdHXABUYUFTXaorBA9g0BOI1FGFM4CMUJIZaixm
V57I7Wom2cJWjW57tBhOKOSQbCboi0YqJmHjGoYYvS71QcvTYIS6Sj3v03tzeax5sX0LXv9GRfCP
VRVTBZ/+rp1tvMKljJ/WAJuaXUnCk2yJUYyOmMU063pKnF15Zs0dIfDJIAwwFugtZ5VGZ5qRRibL
8URso4lWJUdrFhj7Yn/IMj7zeBdRHT6OMsIa6V+2tCBA7DyAxIgyM2iIRy3HM2AZN9ziR1DX1woT
sE3jAEQ2++muVEhLaNY/Yvd3NICkS5ImGn1UEVUqD+4HWcLUJoNjf4XO6SVGUIEO6xHr3Ki8s+tD
C5HBOCcmKpp3LY8hFLjULjVJ133zky2axSrdWlARjEWd13Qz1Ih0hHDviYA5vI6wgNse0L+Qj/fE
RYOi4kKA2zgNfrOUcGV9e70xZMcdCPA6vej6vDUOF8ok69AqmnkpEsZvOkahoXWgmVvSg4HdcfZM
a0UyL4DXWdR428qJO3MyJJ8Kh3Yj6S2RPyDFrwAG9j4iRbkWZGcTh/n/TvT4hux8POSzVuQY9Kry
li6hLp4HPn6b5LfcWi7W762P1ZwNNqGv+3G7eHjpX4UpiMSkxTWV48BfaR7M1S8VGd5LJmsAR76o
uvToVWzKNHR7mOwvnTxHbYmiB60HBMxEA48GbzwlByJ8/gOG3pxuNpQlr1sK/NwbUKeLP/oclO0H
LpC1tZPp1u/UEMKOeajIuNa1mo14b8WJFctfNmYFomZje2GlmWOf/dVfNq491dP+gFUPp56jidpM
HqA1pF+l9gI3H5yCnU4Mb+dU7/d4WXsqst5WGhOBNuJAmcsctzz21g0LNRnN8rqrqzc1CG+KpweJ
/eN2W/r63X3xJvlLgbAWJRdJejSUN4jRXOxtErMEsBdrEIiAQ0zeBm378XKnDV9RfC+6poDWYz5r
shMkWcUt+ApxJXtc8SbhH1OaRVoRX6Dkm7we0DUJcHijPKE9dx94n8qp2ouCN4SAV2cms5lk95iv
whnj/Ebx6ENyclZlS7LMI9NpIF2AyxxUxg2KSTjziAS+ukLQJYEvJ50nz7BLw7X19Og9k6Fnw0wI
6mRumV5KfNl8esvHkTB+Jr41TfsQw6JFXEjqlqefNaO7j81SADDk0C1bIBu+N4Bm2IxQGULBss5A
W8uEuhizwop4pme0JOZ+hJcn7h/n4OVyCMRiAM2qtW3ugddbfql0CXP1ZsyVheVGc4pwW7GzuhTV
dQBEdho9+GeIU7gjl1dN9yCVoShaYMoPq9djSPZFwRq4ssEtR9puKwkFx31GpXKU/a/57y8TYdok
f6q+djBZjRtrv3qZZ4SB+icKWDg5vffI/ybyeSQaXTWy0w5z6yYlDYgDwKsAcg8c3COqDqKap7u/
YrS/lOALejYwKLgUyb2I+it2zWGeezCieyrJ7vwdB/9rXQ7g7BwMFxJQY5uaF/Iy+1ar5+3wbTXL
YNcpfCyrro0xFfgsQtCjUFTjmCCo0FiMptwtStm+KE2ke8XEfmVe+PpVWklvG8u3jCS+uqlIty+N
tPkfWXRWk+aCy6C9jKr4QSrMtcUs12K4Ko55OdIHI3SlJcK6M2QWrd2lKZdX7guT1lWNN22+Yk8N
azCZzn865uokBkdDZyIE5QGxXZnAaxKbRrmHNgxbdvWIRSJy9HvFHW196CDp58fhlZ3je65Cagpf
ZNfhKKjym/RiKwLirIMv7gBSxyp2GShQen3GArJy9oQWJn3F57a6BjlW4cs+5tst2U7U/gXQ00wg
D/LzkIFWqPTKE5IoNW7tUxBGmOlY/yza15A8E8wjlhLRxZ9NnsAKuQiFgde9zBQU+GAK2h33wccQ
LClI8md9W2xAOfFKPKLrO6MYPGpNG6GDbR28hOQIRwngkEuFuQ48To1LlwedFMs62TuGwiYZW77i
ZSAbXANEQIC7QyBXgvAosX37LyeLq0AUywU+L5KptwA0I5FA0+bo9TuQdEKmPS7FFtbwe6hKQrgE
w5WAmq8U5nOjg67iwKygSWmgp+I0m1HhvuGwkVXhV1LFUV8cMF3cLimJDMBS8viV1dXTzSaeNfYV
cY5iWOCJneO41r8=
`pragma protect end_protected
