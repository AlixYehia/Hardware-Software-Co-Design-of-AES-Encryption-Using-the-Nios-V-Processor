// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vSv6O9oGHGZKkDBKQGiEKtNxxQl98s/9E+F9L/12qUDusLwu5TRlRyZfzJjO5cmipPpvAMa41F4B
RFElA8YIbMR8o4K/kpTNMK7sgz9y2yMmTs520rkl3NSWsgECKvyst4lYF2eSAiP4QYrDIx4+u9VR
N5qiqAWd6g9P8E4m009GansTI+EJNfViUDe7A2bX1eviA155GrEts/3PlRHRwVbMq5aE6ABHoz5o
58UVhgpuP39Qc8jYhaXuwhHRaXQMfYfzcRfZEjKoxTJ0PxQP+EQ35iGfIMatRa75N50OzNMLaMRw
buQVdKKM0l1I6WJerhXrhD3jRyXBybZcfBdzow==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6560)
V+9q6+XHvpbCFHjydRXTETacl7limcv0U7eYiBUKAsXBS8mO6cJRDSNw2uBacWRCJIgk71DK+JH9
tZb2cOxG3S4AE74qinWqSnEjZGRhv7N3Wve29h4Ql918CVTlXmpfe/kEFNFtVD4PeYUaiAoENDfg
4RQ0luDe5SAGzKV7v+mDPNZvG0Vn0f60Mdr4HqYvoci5ckZ1MarDlS4HOnGLEChuMxrQOuquEI5H
c6Zv23pdcbM5+jxfFFWXG/R2TZoV50xmqH+dGNrh6Kd+Kv1BOczspAnmgSWEbA1uPfUv/Gu92enq
J2X4uPyksYL7FbUpqzmynW92V+G7/xnEiycrbsl5kTEoQ3ejMfNGoVRfPP1FgBiUotAXDRxsegG2
Nm7c7f+VZrl5bPwoXEREGj6nQ+tZiYVvcKifZr6EA9VgjGfV/ZkB0nrtgYddFiQW0wmJjfgT4Lx5
E0EgRW8dDk8aSppsyE2o1YWRACnoDYdUuTrT2Wl+FIrf4nIMhzBAQ2fVy5MqMLXFMEnFyz04ryfh
yi1wT9+Ga1l1yPnyfHD/e1JbPrh4a7SS2GKkXD3LXHqCB/vrwBNMUPnBhM4LWS2IDdF8KUG5Iw9l
TbHKojm4mfB8Ku0LaNBkuNrpWkp58/nckK6OviyQHyLQKheMgLhI3kvskGXA5kFjJfux7qXy5x9B
suMqtTErPZUkI37pOr8uK+ZKtpP2G+W8JT6P5ltNRWHsOVYsog91qwFvLhWqx2FdM8T/xKgojKtm
ykN5pQ1WbKlVwUtD/qeDpeUnIe1jBR+HDT5w0pSRlB6YcSnEbxc3nr8MKkwb4kIUduxQ3CjQTX7q
sty7oBFgeX8H3qOfM4ItomgVAat09pWi3K8QK2Ac+Bkx8CIk5wpCAPeSDe6yEwkeBh4ewotFT7RT
hFGNKjJBf+s6wG7RYYSFNyJikqxBLJChZjDNMY2VaUHZNXhKxwcgQ3gSmR4LE4AWqdgfG5jKWC8e
aCqJoz0FidYLibFONHtWeM/kiA66PyrqtMBIbJ1nVjreOJJgS7zluvoGDftOICwkZ4epbavn4dYR
HROmiErShAk2SCJgLDwPYwF1ZiBjq2PCP+sA2fiYa5Si7KLocEmAdrfvhJEAOo+c13rGzhvFYr2k
xZVFwtbu4cK7RfkPC+pyzO4e7sHIAvZ3bP7AFifiEHABSMxgXiDXibnItkBkaymklX0+lN63kmFV
TP3R+CZo0y4+YR1808wfo9VQeb+M70ARsOIzjVbqyIPG5ik7ANKs1hzHkbAysdh1xLD3OXzv2tQv
utnuwS9m1CrmpzQSPmpyYZmlcI92WUd9nCikW5BtYCW2ntmHG7kjXXrSTptWYlvJMbazU8EaVivt
hKRaYnJrTVaEIONOjJwopqZqyq0QOqplCn6MVCuQDQlKsvmyICk/iNrWKkm52aGphHrnRgpY5QLF
/IolrvizhcSZwE6+iOlt/h4I43m5DDBvoQWfwRmDwZA3+NhVQTm7mBgv8L5Jt2qADjh0JRjjxF90
53yELVb335aV71I1Kjl9Qq376xtc/erMsZFwWJuwOrZBOh9XyylqoalifadhQH4KEp2yTjeBTvN2
Dq6G6BYhuCpk/BdO8My8z3r2nozR8oKq4HfQAP6ntqUURrh3VIF6I8gi65T+1AYMw0IpKKbVj4S6
DLTQuBbAnQxDf6U4hGKIzss+Ezj84gex2Nmi1NidjfmufRcuIa4xiAqhd6X4iLPQr9MUOTdkVewi
SVJW6+arEO087I9dSB5bi9Yr/lUjGwZ/ORmg1mOb5WIKSFUdvL0i3alKBfvZt4S9t9z12TbQbNo4
VKaEDdgKDKOesu/yBGngt2pzqzUfOBpY8Xv9ASyBQPiari7ieXbo+czQuKw6FkyfTJz3/0jFkihf
YWDaf/6CvZFW2NL3/1wRe2Tegu2B+FgyC+IzYhex9YmnTeTL5G7jfj9dvWCovTmiIWLeqgoTFA0Y
5TaWyA7C3I06zN1OYoYoP84sZsUozXkzaSmRoYxFxpaNo4BHbGrHn8ImofMzSEF6IKScz5LjpE/g
M/XIdvI3e50F4iYpJvn6QLsHWe8zr6YmmyFLmXErTAlpJ51NcJ4JBRD5sg1rPGKg5BBMWCSuelPJ
ymDWMQP3BjusBeuHshPu+asoSeWIoKvQTN8597gSsgGMvWq2FqpkJlgWPRZMHBF8oGr1W3u38rcA
tUveChidR9r+7+XacXnC7fQFFuXq4ZgyuNc5xwyId4y+4DJKLIx47h8OVQ4IBe2LB/DhlIY+DOO6
uR1ij1qC2+MlKNdg15BAmzZexicDN29qJ2m0z32IpC5ZdBMojMUqU53BLBfWfHn/3lgpuwE6xmfT
a0HP+xmYu0PXEcGs+RufkRk56I1WCTNvHMjQHzGRa6NxtS1ts6YhxOTY97UAGqf6Jt94weu2LwWh
xd61VEY3pfWUDDciNLgCthPzm1j3qSrVDmBlcofaRlfcP9EfpJ+9iDnDs1sC2nnmEhAIFFy0t2qY
1yO1rF5sIJOFaxEXyqWD8iVcp7Y1jdriGOnG6mCxrSF2SXC6Z7kT8gYu/tpMVWapuar6SD2p0D3c
hjf5knMpT0i8iu1zyTrRQR7o++kOk3+DdfblIlbRcar952PnLJbIeb8Btmm3wH7c2uzSiqKnGhwM
qHh1VBt3wlPdIvQjKLtecPs/o6NkJQnVctZbW9pFsTskjZ/ZFQKeheHW1PNoIVlOJ7wnM7kTQPUv
+W1S6tUD/kdl4ap9xrlf+rJ8fRnd3SEda4XJrh6YegPWugcV9N2Y999j7AFwi+jRIeKEqSnkkyE2
NccZYpUkSgESaG+dPCFx75+f6IgxZh4I+87OQfDRpQEIJPhO5CL+7sOSPSScLQYOCDg1mPlX/5DY
jxVc9OQsXyUsaLv32Gvj8FmDOfJfxBVe/8fzGjonLz2YtRUjcaQ4svCiBYV+Y6qx3Vq6x0XoAYvi
6yrbkhWS2EzKkNkSsOf4pwpHa14l/Glthi0KmovfCO4I9TvUaaO82EUg/Nnc5GyqTkEA1Xl1Z2Fu
5n7OcNlIup/vgahyXSnlmYFQy3JUUtErKn19OD6lvA/Ei2bQxFGOOP0aork45g1/xZkPmNFweV7l
qRs7zw4bLaMgkDl5nV3Br81lqHdf7PzqAaaOMo/CN09Sb8PtbfgcpvA2Z3AKtAKNzrNbcoocmmiE
XvQZ5bjZUfGsKscTFTNVk5DVSZZUpr4F+LvHFcGOnsoD9JDx639EbqwimmEq0LnUUbRmIAbXgfp7
uNY7U70EVNQMBid1GXjAfxU6vAxF3dubaU43Fb1oItFjn/onbz/uv9PoWv6DUXGdyc7ypgQTBT0V
WzVopKSrBurZ3niNremOyroGmKsYKHV6FSwXXU5mQ0Pd8YVglnjnB8sPWSZwrDWu3ZN73gImie8R
2X63lIWwTZSgQfzG/Wdipff/QH4yt+YmPPGctheRPkOOt9cHVTRgUWTd26ujGVtv57xBMK+NTBb7
VqJDEpZPqZv80sP/DWMMnoHSYOGuXsHSZy+22qpolT00UN9P8gBDwzp98q7vNJKk784Ijk5by0sl
7icVnWyjFqZowdL69rJxLvm4kcnFXZ1SiZNu7vkT6sdvwY8JKJt/gWe86jOahhwzG1RTdK3wKi6X
DfeJsEQJMp7SvksZNoFZcnF7A1O2SfRkSziE6dNCxh6X1ZnpgrEm+77l0G5w/Ki5HrJc/O2eytSR
hwOq3WgXwIoPN3MJCdzL64bKYaQ3B+8BcT/4l98wr1GQGAiZr0QChotPSGkR9nvawmXZI5b0+0oB
m78D0e12gm4Gm93HA4OyiqSTEXWSQdbHdm20sysbFON/GLz1rhJ70/DP/cEc0l6nK+j3Xi7s6Im0
39smUYlkd2UMHgmgS6bRcDgeDm3yjeFEWQOdF/dDOji8cfC3PORdNrfgqjHhBRVIpaXUQ9zaTbyP
V1h4Gm5sfsw0srBDsCXhZ9LBuxjJGw5nkLpKp//61KQ//xvgedIdU1j7Dsk7hDaLv8o0eoI2VGaF
r7WGv+rrggD6AIPIcTmctR2Q6wOGAZu2hAWF+HLvzhswCJePeuhdAFqN0BVNmW+9GVmq2JLqExD0
UhDAbetAFxPaSLFZa42PBUsVlUWxsjojrpYQDeSc5f3isTtw8zrUoXxwle+PL3LCBIwhpjICiaNa
E04h9lz/4AKPpfDTWzcgwxwudBS22FClFNBH015fyJsP8C/48CyCese+hzb3+jRIiMbfVfrLJrkd
6KQh9uKQb7gbgyiBjG/0aITpOtFPSZA1sab5nEu7HN29+9Ew2rHySp7Z+8ZkuxHOwxZqkn8k+Juu
UbwGJ+hUzJsHHXUPDM9B7IE8sqkv9H/dDNMb4t26J3VwSBHljZdVqtBjPYqQDtHWcZ1LT5SA3ibJ
Vlxq7LAzA3mcEWZuHuq14ErraSI/vogW+trBgszh+MvHdKidp0tx9lURLuk3BaDZjFFnW4+hZv+G
a4g7YY+wIcoIhJqdFYY/VSkZfASyBgSMeTZp4FPG1dkcJpPX5fMYt+FbQD3k7RQDlJCrtK1R/17T
obP8YWBBTrTTlag6bKbQGOdmPe/20naAvynbTLyXG0M/u2G5tWlJ86DbBd8g1RmRh80/91H1s62e
9vckf/Z45mqx5krd2PqXPmYmpbJn0oa916fSgCgsSfq6DtD7XxKH0jmWvIuYfZHwN4VJcCvchsob
PhBU5IvOBKlRgkWjK6lvCrV29CxBCDv9F95tezpV9Ile8NgT6rhkf3V+vbaY84lzeRmZgDLONtI5
8pHvsJqS6K05L2tT8nrAaDHZQl6hPxuxtBIKX0f3BAeTZIOTf4Z3ylGkWpPdcCVDKs8Ij2YcbaxQ
PQJoDE0aKgXdGsz90DE1ScDABfoU6ycgqd/L8vMHc6xZ9SZF9HkXC2dCb3bn9OHwUWrs4lZzGCUY
WsxOcL4dRbzWeAaEhY7PVVRFxMbZ99cd30YPX3Ghnvud8gGcuU37dbzdhI4DRMPC0F3DUhy8GoWe
x6hf5ms68kgkaQYQB5JZALwBzA7MuMsN/tLW8flZIajxMC6+rs2e1V5d4gDTT7vELTm4xEZs8NdF
8ajToMqYlLeyEn/00Fkn9Oj3dlvt1I+xXwoQdjd4pX4hFxIPFX2nXgLi53V9fLfPAkiZCD13g9Zs
kS40XutHuZdvcUckyckRQMiY81O8LrL8/CvouljJpf0AdODql9CX/INZ5QVrGS3BlCAT8C5DcFzP
CkRFoHA45ElQLRNCLJgtkL0nFNfyxdMmyB58Sn1NeilwVeYoj0ZWaibXmuv8DjgWoJ7IZGlisOwK
EXtLft0xcKXiXaAchjt8xtNczcQopb+LFRiEHJYxn0/oljJrWFnRwWZ2bd4VSs9ktY/3SlczsSAf
YFPO95mxAsaXny8JA8EpMG2H8Cdc6feA9gffHSsABXSA5xC4xbivHwoEhbDQjUMDMyzwbXwYngYc
ujzCpZYe7K9QvcXfuaqTbDdJbtt4ObRIg341wgfR9kg7CUznyPm3tshWOtx3FmEbqGD/QFrihdoz
wA5UVVZ0wK/h2jptDLsHg9YEYu+WnCBuIeTV2XubJUCvZ/C3GkxD2edRIcmJm5IJ6AENfvC5rql5
a/ZiMVTcnNtmJ1kBZzbBofpK0oXAkRZnaxVdTibZa8rXIi5jrVWYyo56P5WcITHUSO1pgHoQbX1L
MNFGGjV/pM2F3JN7xwhQUjGRDeAZ3Z9qLasFH65EbnNSxJnGzfY7H5rX0dToRpwmjC5FttxbrIHc
kVJ0M0H0LsTjNViwcBNi40pC/cBHk22jyT8YS8IbEENBBvWWYhslaXZDPcpMSEZoD1WRbGn/jtv0
g1K+CdjuS7dh78QXo+mk4kUvEtgsR41A+k+bCtsEdh1/5RHQKhyzFeCFCzoiBUBNen/s4WDx+Si9
EkoajKZHVmWcGo+LXzjot8vTKysJii2zLN171dDjKce5bG7TSWLzo05Q80chIg9GQJnaJXNxB7yc
QTGIYEZ3QMo9gjpPjhKhoQszdl51bKVlAee0dQ1qSS0QAXhwnzIrRpliHtQ0wMm9aweucGSk6024
hrp/t7Gw4IZ0yfpZdArLlwjGZZ3DshHwRV17EWeG2yRMNbj/JPK68gCYqRF4TM6+fWl2xfNiy/zv
bkfuQ/BvTET+uy6RGHheZaTQSiKVFB20fyIQbc6bBzwssYvdNY3mFdg3Ni08p4C/8702V4HPkIHt
ghaFlPPDTmfGrVqyvHAyj7gmnk2TlXUSdSPnKKgq46/9yKcN1hZglp/ncbxtSghr7o28n764lOhx
zgsYE4QOlyW+WltCw98WlGeaS4AWBTuDyG0e8nSKLViCLeRipagDwGww6kxtOqr/zxo5+yiXpapi
mbEQ1RmuBs+aS/e7cMjnM2F56t5pE2mc63rYev0P1zmkY4Ak0zgRfxhHFSSyhx4LwosBjxerkA/I
sgpBlXFj4QzYOtT+UQxamEsECQKkB4pvMmr9/me1HO/FosSxADx2zoihooFSKEHg6/TNNm3EQ3Ld
qMBuGZasNOrhwGbthWLigP3W/9b2uoSQy5ctJ03LX/A77LtpQ3SBfthqyMzHq1Z/0dxhfFzf3gek
AbtEleAORT27aOUEgEX/PAN1Uo6YI8cklPqjyR55rYond/Xn6igpWu4qkScyrmSSPb5PlOVxWH2P
93FxEiFyCbj3sUUqatgRi4Dx9vU9WBnUziYT/NhHH0qTkKwowcn86BKYFCgHd+y3iCp1lQm1qvSk
mYXSWw3g8xvgFnXaroc4VbhBoSpE9MxxCYWKM7MJHIBPY5q4pZePP20eDnWTGTYyXhBDsPSymdNc
3tz9RYLn9z734nNuX7spqt6+uzsisM+jWUoujXCJm0PE6Kq3951YUX1jCTTO4gdTQg7sm5s5yAwU
7Q1axrHu2w33408oAhLMEjzuLNBtWi7gs6iWnkj2mBjDhuIVHDZg+4/TJH5Zvh+OXby+5gM2srLN
yvoEqGVHfI5G+TTb4j3GzPTg1urYRNoL8RMF5SgtCljuzPxakUmbqkca/ADwDyn9Bm9mSLKDH8dw
0Td/8YsrMw6kkijOzarxVcWX2igqEV0f8NqAwqskxA1dG7mcy0BiZbeo2Exd7171MhTohn7GWcOS
vkMXzMDKt2TXoE9XWsT7T9wTlC2cXlgPoUvMyoSA1oMBGASpHnJ+iRfKnZj/shoC+E7fhT3NSu2y
Rdi21jMFzqopHMswDX6oUQyu7DCtm9GDvSXpjRzYbQXYIA9xoPQmjZ9nVYry4+0K7YXu23+PZmN5
BjBo7iceZt7eM80OG7ecfgYw/6P84p4cGulMr7pUbeV69FgGToMMT+StDRlpIvh54QQopuVUwJmV
MNpIj+3MHGkCFwE+i2nq6BfuX1mVtzYfDro8+7cWWaTB7Tax6gCOnPxA2ZBJu1XENLcsRUKV8lTu
KLvXcQ3C/422SHAltnrk9zUwuYo6AV3DOlY6khEKguKv+Ai5OjQit2qKWZM7tlT1Yzjsf3TL4gBU
9yn4mnJXeyehNgdEWHmfOqItt0kNb/F2/DXJ04WwMa/blSFhUcjAy3Lzjb4FjfyGEPlc7VLEPkPB
SeoyvMPZoAT5kxpxb0p4nTP74KglhCVB2mO7CKlxkk5GlajM9loaZJcpdF8sVgXTRLzNcGfHCFNf
vovaU/3FBwccs4VHr1zMHJ8q/TUKyXxDZSEvIDQjRHXH2jFBfW00nogQBsD9aUQR3ECWr7uLsDOK
CypSavRGKL79PAGLJHqCxydkBtcpDx03FrEf4R3hk9GyV/p+FTajj7M0jyezJF+vqm2gIs+WwUIf
C6Uf04wdLyqZU3gRGWIj2cbOVh7ZtJprWLtErkQOF2bdc/zJMUXDaUDijRb8aAHrHcRhB2WKFsML
oTCkIzeSewD7GnKTN6AfPgKGNxACroX7gb5wMFUAXWskb/RBtSKPQpCMGdJ64/C0c834Fo4gzyVI
l2BnVNlfwAgxK/1pYLoH0mVZUcBtMvs6nnr2qyHO87LBz1hramk9tqmJe/k1huorlrSCQdZAut/6
JGglfJq5AvJAUxzgOkeD6TWkHRYnPqGomBXpVpjRRrLfqiRTS1kglHrMMJaDs88LEi/5Csg5hWzB
NwHfP3ngNTO1JPnNhhmSwHmEEM38iJei3686QFx+iiB7OoDmUoVdhza2AX8s/yOo9c/6RH/+CgCC
/uhvU1qZS3Bu/GH2wNri6qruhQvNdtry99pOFY1/FhpyoqnbRxojN9stpexzCBw8j9IrIQnqjOIp
HrOsJ382VJcHtpZBg/bDRWFAdqASMwsmtXOsUFoO3X5+OSaVvtPG8wwXkJmkWevl3KseV9nuQONi
hf/RoYaUyGUOmuyoOsnANc2bMk4KCA4xmyUHHTf2fDcxrvlvU4bftW6Zn+RDKQf17lOskHjc9J+7
OR8KTS8fpAwRiYa+Zw4VLTRTmX2NNLyGmQN9rRekntEWCOKep7AZZHx7dNgrC6h0RbwrR4JZTpgi
dmaE1cQ7boVCXDgzhMesoaCRpL831QMf0nUR+gSmmoVUjuZ5bD3nKGZPiZMS3olcGw2PExYSW7jX
68M4VI4mScGJVcW+TNTwPTYneRj0t80CsoZ5A5N9ys3H4pRSUpjy1oJMQ64YUktwwN68f+hXhJy8
PNCeg/Ui1wHAIFtVZGJV27eQj3xic5HBMt2cwW4bitVI2t+RXJ8nrxh9yZvvZ5bwAdVCG0xX6jPc
dU2NWB8=
`pragma protect end_protected
