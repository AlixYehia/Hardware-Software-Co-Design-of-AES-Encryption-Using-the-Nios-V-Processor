// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
xlS02pigoiiLsgMplEsX1WP5UiZzVNJ00Bml+d5gRaPRftODNczC2dKrlDiGbmmWLbw+pZ3B2rmK
ubfBksNQkXTk0r0GOqO4MewImDMU33oL8jK4kqDGRBuw1gkTskRWYtc3pYCVCDVi0PK7411Eynum
6mbod6y2jEBiWTaeY7+39Wx95vcXfppvA32Qsty7g3H4cCWawye48PqeRYKWk5D2Ah7r55CBBhXq
Trr3R0uOEPWQZZq8iCg9QkVwxqbEp4Ew0HBDihiwDEV8jOCRIU0MIYInwhNG3P7S/h/41AW+hTR9
jFknUY8eC3UcM+YhMjd+Rheynz2nnejKy7HWaA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11184)
v+QXrcT0I2ogpRIzdzGJh7aQAX8Ch5N0btiuGzSJdtOq25z0s8tIN0umXuCnHiPAB3Exy+dQrLbS
WObd05bJ2D57mlVomrBGelG5f8NhefJfUuRpx9m3OLtZvhS97Lzh9f7LUZl7YDw+/63rgL8nGp30
C2/R7bSEmTB5sKH2gUDiq0YOnafG2OU1TwkDtw6SDRFSumj59VtpDEPpWxLSIW7Kw/P7PuRcc7Ha
Af+crJomsaf2lVPookJmNxlRcDGaFyugoAwNdE5TA+FxGbeDrNIY6n39EstQisVyjgu5qrssKu2b
s4paRmrW6Cv4INjhRxhr3SVrmMJrtGAB+POyPE1eX88YS3RDPKOk66XeZiAHc0TNQxKAw5bQ8kpP
FwTRedngwidvCTZm9w5Bm+nlG9aLCNpg4Y3Y2NwyF/iMUeS9SdZVfHlHQhmEqPmEJI47NIq9OWLj
fG2BdzZVOGc5cmz2OrIPgMu0E2LK7FU0o8r1+Z+e+UthfPK6MKeb1uYz+0kWNEfcFw7IspXHPinu
Hew498XJ3oTxTI65dRD2NOad0oy5T83QWwUc4DFv2Rk5B/ZPand1QLO6alBVjEcqZZxCIv6YSGwy
zEm624pMeTuJtVLEg/Zmq+BqRZTnRe/Tiyk2b61Ndug2aSRa+HTWsIWuL3ah7KWQ1u3kpxwNALKf
3K6yj9ahrE0wn8rIbIjLxTxOYUVhTi8NCZ5/l3Bu4zJuzLmpm59DgZDvpRr/iucqzaOkjgn9ZfZ2
+DCE6+y1rj+USiCn0yraiWGnMxX/5I5BY1d3MCG6hTrpRYk9wOvPQJXuuVgDcyG7AJjS/yZ2FW1f
hiUpfav4WgIESFh/XEG0dlAoNAHvg+ssCZax4gMJSBTIQ4ObHRK+TVGWVtTMF2o9tmj0EAjye58H
6nRFblofTiB6Lp8PTpQx98hHXpBUdAqBkC7a9darrSt4B+6lgQvRa755iM8cV685Yf7kE4jfInyL
4GfQCZkQsV9jfu5NWyCcCddpKyBNqxbzsU9HeP4R3ZRhW/Zlgy6/HOKcBxXHKbxqOuXs7BYgvfww
PqRYE77nq8Ll7pfaZd+x/aZMWAcMP3LZEh6M26mIZQB5ads6ojrbPdXz7e/510eh4bNby+CgLphj
Txi9cUgHJGeF5f/FCbphBlKCSK6894o/Aluu+wTYE6Ve/xMEUWPSZyizEkfiSA2oSUzP0OOXQc31
yU3FH/FQmC/53BMUVx5YU0d1PyQynU7Gjuea0CT4Ak5EyP/0EOH/1BnXtbYAjSprFQogxXdRW//X
6k3fAg9WYJNKvhkOW9x34sKfn3/XwS0eyVPSjvMXKwDpNwh5rns/fqmmYzJInKd3LOrm5dMwYGs1
6gXZgJeCdOzCazsy5p3v5gc98db5x5hE309gxj7IbyE8SeunobczmC+A9UaAeL//Is0u+rdU9Qti
U5AQ3pLiMeFIOiMsd/q8GBBx7vGsM9drubuNbvSgAx+rD++uHm6nzS09wS0n+4czpckWjqqUPIjG
W1Vji8GJpUhSsjXUPFf1tsoC3FQ8/bj6KZJC0ZJLzfXHdxQT5cbnm4BRZAYECBlN7tbHa2E4fmnx
cBrqRdfKH3w7ILqgRYv9OBlUOhskyfRYsNIeAY8/b8obRO49dhUecoWlgnBkAItXrii3fEa/k+zj
H0sADPh4k2gm3TGL5oiqsFe3AC4DfDMdOCZolY5PQyrqaI5D7sn1gDCffTnYri1XQLZUunJ9VJKR
9705kd3PQFNAZtaA/65GWOzblAZ694FEDjn9ZKs1aoEt4CzGMuKujum1fqA2+glhmDxpQzx3dOoq
HI9BGxgNBLExOihehfDMoiChk2A2/0cfBGnGOqxZ3GvOSgvefOtO+2b64hkVDglccjfFfmWyQ0av
ZCzZQZGf/HyDwYMcsx6IYSwV1vKOJOYLcgZRwthJtGNRYzROwOPBRE45YcfU75Z5k8Bbt4tIJqH1
PTFmO99yQiDnA1h3E7M0OdBNbbL56UABBjB0lXVVTLJJHq1NdvtAt/KzbuNqiC5FFMvpsqGerRB+
s1/EIod3DNEI9+mqgynLB7zCr+EVkCfor3ITey5eAGcBDEZkMZuot2SgckvvChoxrCWk1B4MuKLv
A1QHCTEbabB6cxd9ikhHCzYCtLez9KJywCbTf+dUX2DZSlQ737LT75KLF8+ssbfyKI5DHb1J3c6S
jUovWSR0ygsH+jVloyS/2IQmegbHxv3+2AIFhgYJ0ZFCN50Ipdgb0TnFsl7cqXHFTcD1GuMHVVE8
TfyADrgTfoEOeaQ2cZvKZ+mtMjmh9gifpnADVivgFNpUhCZz+iFSwWbYptp96ijazOFr5fxc70Li
ipCunvKIvzryZ42gPVrVkeyMloee+RvTtkeKBoAw0vcR6u/3Viqg9opN570yFpi8b9QyoJwlhoWi
URZK/V7vZ1NTSUo1NAVe0etlRWsSwa4ilyWiSBlsn3PinXVg71tbzO1zj3gq6+CL/fO3tOSk7Ecq
1wcLD5pZs+K6LmhkTinpBhP0Sd9KN9zSMFo4H2B3H7poyOWkEk4mFIgiAdE1In+kiv80hi1Th5cl
8ZNEpwuL91Z2YSOXfEkEVhq10oZYTGgK+kDa/zXBbZm6PNUHTrNET9jQ+LoYbfHfY32CrPblaKZp
Agk+vuxuVjdiapaS2cczTebPmqTc2l3IJrTikK9NkraI705UJzFUsUMQoFk5Exz96OfVF6TsQcmG
f2v4U+H4W06zzUdp/g1MeyNqt+OL+TFPQOL652Rt3HLazz0L3TMPFelKyvXLGJJopAAyQG0q1WPO
pyaZJ3pqU2UcnjWrn27Ck+wqSNMJvnRhOy43IDOSntbFy8qiZuY9+Uuh08LxnkGWkbO8i0bOVDco
W6kUt4fybIhdgOYK9Bqo/LSYeAk06PfUtFagOe0aAhYKUBfODXmXVlYQ23EGJGqhYVtFaXCD/hG3
XOZbwKOqYymecSCaxWvZAKtCpKYRXCkru4gPGSg+Nr3dOHFdILWjIsAO9itTOAAL3BlB3K62cRIG
ANNm83Ma4GLlsLHouksNUwRyzMfE0Z4ZVfywHrk4E3clXE7LNvValUlRp0yAtkoJpZnoyeCGQTyl
iKGMM2faMlUD8VbfEUYBCAYEi1Wz2DwtkHTI4pS0ta7azfKlyMODEbV89hhqoBDcd/bzOuEK+88A
oeCXNxTNkLe9uOsaqDxBZBomlWSwPrYCWeYIN7xh0sKb8rn0GaLI01LyhJ6mLDpvMSdCxWGi8AgY
+Dp3ga2lnMxcGRIU0zQok1WBelObTFDvGfbhD9SlHjTqM4cx3IGQ7bDaziIJARw57wpRrbvr0OKd
sw5WZv8yPqUNZazhwaizUx72kkbZaVVSdX1DaBF/Bz9GQmxabRdOKP71ECUkBUDJ1/GbhAENuMCB
j8xroA3+5KyjvPGSeuR02ltoWBxh0c2VTwvKXq1XKyHlbIiqZ2Sv1OWGShz43iB27Q6dCfT0UDQQ
hK/vO7/VkglpBaVwCnNGpCKst/+QnJMOvYGQwJrdYpjMukGUyN1Yb9J4K+Nwd1AOojg2U+MTliIo
NcZB0pEkJuMbnj9maYkDI/Hm/CPy2lMqVJ5azOw9oggnMmmRrO9QDTS+2K5ft8OBIYv/pmiDOTwd
F7aRTidul/SnbMok2/vH2RoRBm3tTYKuYLEk6aUwaF97nhh9z0nlaFTnOEGgCU25rbfLNtZwU0nA
Uv0s6lF6WiOV6ClMt1SwURCyUuLwkrk2vJgYUMcsl55NiN1ILOVVED3Hjq3DagDdYrfSs9kwPHmx
XQIHQnJIZIiZnR3mU22+7+NTvfYhwD6iKlsI/opyK/iOPuMy2orfoN6d5XZP8i7cgocw/gnCuf+L
f2desVl/sHKzv/Ov8xCSaqXEqpHLsPR3dGWYn+8DNNwuxjJc7DDnJqpq1HtLgOn+3wFdSHB+Rwhk
xCnUJdomCeyeQjPVEESAOSwmEe3M67O3WeK+8L4GzQVlaj7SwK0h8G7EwhAinpZ5MV4DgUanvieE
Sylnuus4cESrNPh0xErG8J3EYGmRXOsB6+rOWiK+T0UBu0DPSsfB1JoISA5BfUcZrfZxlZ5kRrcW
BRRotj0+epUJTQyzminupKfFcNTRoKFHYqsfuiI9tC+Z9WLbgZKvLzB8SD7gCXCrh/ztfE1tkYwn
dVFP6B32iNneUwRFeyrY2Ojyf8XSNFaLzrCEjuUA/RB+aMTpE8iOoU4hCPg6R1uffFAkLMesUyuH
xJBPuTprBGDLgyzjFtnSRNMC0W9URi/P3uHXnn47vs8Jf/1RTJKUniUmLr1K3fBbpzkI9NYCxCcc
g+nI3U5CoDozOos+Is3vTZIHmBA75eDxUrxwEeXvBJSo9QzoDau35TkkkggXfWhtcAX/ObokrYX2
rLvlchU7Gos2VKqXNFzBNSJO4X6SZ5zbI8x6BjpDpZ8UfsWdlPsDw1a5SmxDCArdpiF8lFiwm8gO
P27oNZcjUGxLrbIrpDk7GIT2+xlZsAkr0T/CV86dFwRbkStbNkhbFcuzv+O8ZxQ51l6ZhWFF9WnF
9XAeo7oomY/I6mnzzusx8nbs2nMzCrlJXh0fBQxvNo9UyeHWYndFOhSY8EQc9sBStmcCrzqjY29I
3rvUIDXsfETSDvP6G3et41AfNesocWDgRIwCIP8izBo+RD6SLBV830c20/8H7q1nNbTHbNcC/M0M
Y/g64qdHS86JnHAVPRABMubNlrLl/v305JREX1/Qzdutm7g88h20Yy+kc7MCtGWpuZRRNrSLDWF5
HXtSUVDkT7/BHuPbZVQIMIXLjbYYMEWKizWZ6whflzsLqA5OcJ7AYQRseu+yvghIXBHiNdIomQgL
QFOCsLcyN/jMyIe1LT2bKsGQOH+UBb78rXc1edhXEaDWdg2rmwr7Bp9FNYj0mH2z23/Vh4M6DfOf
PMqqhv9525k9huw1YRfxDmn7vXq4UJYX7ORh9c0Pcpuz/TzwemMbIJht4NHt+yPW1E944Lo89dmw
fAwgkTPUR87FF+hvMzM0I1HKA5RPhidJxDXom0sIGRC+sO73/K44e13KIV48ztxON+Pc5tSs6JOx
rFIjIBztW/43aNrxznAANdo3NSwrTPf/KbhO9qF71mJq1ghjKylCae16x6W9pLqWd247UzPFEIhD
0BDoCGpD59GQykVULNLR3eKKIZSquztgLOoalT12rdK4Z6BBPiUauAikagEjyBJaAqRJdl3bQoG2
QM7nZr4xDMeEKaljOo778ItiBvy9jo+8Q2V1S/4yEJQB5Btl65s4lGFmLE27e4k0AbY2+buGXqgA
eN8yTzg+yMYLMjXREcNlvWZsS/87g7ci0iinPATPUvLYhdoqnttZRRycF7Bo/bz41lZ+COkDFJYi
nwHdxW6ww7Vu9ESJqfMgeZFzBUHLvEqN+RDD/TM47vwWCyLtk9gdQmlHyU6U6y7b1D+38f+ZwSKu
lNyCFGUqRi9zWdO/WBcNMITxHCgiwzzviSLJqyYHbgrDavPbz5UsEPGoS+duyqh+v3pl4bokZWVX
RvLfwN0PaX0t7RJLtiIXE9he252GG1OQ8xH9k4ZVl5QEOv4dWm+arg3oTESuW2UKoNoMx9MbQz+o
97nkY1yftl8VzmXJbb+h7D6E5pdorILKS7qnrL29Sp85FbC4RIwBbYVbgrTXlLjw414n4MZ8vZyF
isuZ9+q94vRwcLxrL2WVgjDAJRazpOESSNMXsRImSMjVoJ29NrFMAaBjy0xZ8/NKg1VmNhPxobvu
LbiMnp1woP2N7e8e+iWyPAuE7ljmyUJvIC3ogUysRfckbw8JrTC6EmTV5TVcAXlIaimE52G0djKu
obBkkaliIdQEdsP1TpFIhFUaery+xo4cRUvGfCu0DXZ7mo4Zz/hPvZHXdaLlcxZ/n8DyB/IYeyd6
heP1jQHxSBymeKUWoyHXZbegKI+v0KlGQx8cxev9vmTwRdALg0n15I+i2SHV7TBWDhIyP+66v8wg
pEbZ519wlcmvSVRcDTn9TPv48FQmsjZAoNPD5B+oS4qMUosM8dutXQ5Gd0bYfXEwxJIFq8y+HLC9
1xJqtHHKsQoVWjOMAoyup2cghA0GlRRvJjTheTpQ1klvU98T9V2i0JYWAEiVw+C/Ipw7olYlhHzs
kBYRCLHH+UcDI9QJMXEiaVbjy4l7ZPqIVvCO/5GG6a2a7kWmhvZP8ujir9tSV/fPL4hxtw6csnTB
L8TFcx3bIy7AqZQHGGIv70B+oEcCSHhx73FGUWIxncE6RhTfVy+B1Fy+BQbGDguiB9bKkeqr2GOY
E6Tm5EAjC5bSzly50YHAQjQTZnSlH8nbaMZ6TWLS0xsrTz8CMsTzFpVU6rARbiNdwAge9E7mZqzN
j/15mTheZBBw3sFECfuQcQJLy3AUIDTZdjfEz8Ij9To9HpNQHD5hVAwtLqHSiTroZ/lhM2m3Yztx
IdmMMijW/xbOxDVHR2bWWJywGvZcDoTnvv9Nyy3Ze1vB1MZJ3HyEMMUe744WdLqAPPGctUKZgeHx
S3cJEPQrcg9nUqZtoAEOhYnbV9bcKtTSehTTona4TshKDmSrx7ELHRzm7mo2ZpMeBVmKeh7bZ0FB
Dwsca8glRbnAZVW0rTF4wzVmfIhtkcBLDS+tmV5Uu6qSbDuaHQZWegoso1TU6PNNiJEVdy/GyABH
+oqHK2/Th1fwbLw2b1h8eWSiMpMEmrKwWUPesaO892E/JMh9mccW+BiUkW2l4zmgSpOHw5/6ioDa
cXynSXNVj1EXX69oSOAhS9zuKsr0bpVOqOccJCLgBZItAsV0sdKur3NSEdBzKK6+2cnpxgJj6Qol
5sRbsuvhQxkrnhmXvtXjZg5GRnWWvIcWe8nuFDHXIXbJ4fgATstn0L/eS2tHzMcWXB28YNpfzPWd
qB31PVn6aVEdOnkQlcYGHi6XmhthTShiJydhV+kUgvRdHawUrkqI3jRofmD5juQpDq8cwK4j9lPF
ef8P8vmOIVvLug+cGYxN/m7Cr8H31QciIxpMvbkNScWgoidRd3gENFGJ0KGSyPdGNYgKQZZhuWrF
mRclDRzV/taUmrpshBnD23vecDt6OyLh2FM+vl+mBL7XkgiAr/wb7vPBM7dBeD+OY+am0P1rPF0v
9GCNwRVDoeIljDTVC/WdyIUTFonN5rGoqZGTRBRKgErufqPB030P1ZIppkGqthTN6q77dtdOs1X/
7Rv4f/QHzgQUhYhQrsNR9ndfHFs3/txNwoufsymZ2zAwGiY2XSRFJ+BU9dZQG+hVygdq+nflA2tc
YgG04y6s8asYJbPC+BwATjpb5gOIzHQX1AT50KMyeXdtlRoV7/BY7vS+pHDSWI+qT+Tc5xuJ7i+N
cb7lcDX7+7zb7cQQ7mmucTPDt0zEKbjDDR+6Ij9mJPwD1+r7Wi5ISju0b9gp7h3tI5ME1DQU9yPA
0ZRCxQTdh8cnOqCWnivZiim1KhCTVuDby+E5o+QLRkxfa4IWoVScQg+OCtNgO51HOyivv7a0c+yb
Dv9G+MzGP8ktPYVscyVbVZJmee7RQx0tPFeyanORGTNCmrJTGpMndCnYOj545tDLeHh+5oo/2VaE
GRLjo4hh87tVcqSL2M0eJnrbUOq4yikVBAFkw8FY/uUSfh+WygwnzsTQNAOACXRjI6fEDh/LC8jy
w7q+5PB+YXSAL5c0IAl0m6wZ4J/9RrRMh96Orb4I1Z8N0pKV5U6eFKfzAPhy0iheGhnieQ5yZpqY
RKZC7gA5AsxEu98Ax0Rfl+79MvuWe0SrzuBcV+n+m5ZagHNVgZS2qYRaym9qKyd7oshM0qAJgUTJ
E1CYOUYTFarqDCLzGQt4nlbQHO/6aeN2WAZW343j9VDuf+Y+ta01Isb211bEIXyLkcN2ZKLEfwrA
rjaV2Rxgi5X4RG/luuCG8z2hA2FE+wnaxPEm1YBtwaxhJgCKketLaKpZQoqEuC5ZwseziNgN/+/n
gxZp2CD0obpeFFm5QzPXg9iw13rtlyz6aoixx4ALCJLme6E1DV9CVIbGD3BYwFI0poNfbQ7ZtnFr
UxDNUGMVp6/n7GQqTyhA2M0GbQQVlKghN3gKAt4diNZMAWzFyMONcsuzsPj6LU+iuBoYVVbYkdCI
s7lapyiIesWp6ewhV1Fn4XcX0K1By+bdRqPNCSayDptHEccWsSyu6TfyiuzHEvzliWa2EsMJUCvF
2tt+BlrZc2zB5PbM9sNttMDlm/59mG4bqK6ppd3b6GGsm/6h9SPduqyQ1QK/nYgOTMyux+nWkroV
CxQKY6qR8vUw6gGOgPgoQJpQmMQbuPutkDmSo2zvG3ojd1Mny6FSglysU40NEdyBplooxi5mYr89
kzl4dpgsAMNx1D3GD0iMRBO00+zyjFg/iTyocxckRjyxTI5MIQgFjv3s8F9gbf5hXOMHxRj9IFR6
OkoOU4Ym9+npGfjkpkpTUFZZgr96iATQCHV61zotRjeUHAHCpFPJ7tqJVpNnkLupW5J/XQXvRmAk
tCeL+OhiQ386ar8SzYxQiFEG/DHq3l/PbIMHu4gqX5nLK13XY3IFA3RFZS/wUc/2q8nvAkg4PwRc
A3OE+k5L+eTcG2GuTFt2tM09GdgVche0fEOh3M4LiEIX8/8eJ0jLubhU0VuHXcO0jMzDjKIsBjyG
VQtNlkRRGeVIxpo7GXs+55ImPLvNIxNwYDcQlHuoNJcfydRbOlb5VABWLC8ZAkxN9b86qffPuAo2
Ec46EEpMUFjNFSLEJrRRMR8tW10a9AcCJrBEM7Q+paXiZDRE4PooqAWvAp+teTg7ybhUcv45stQP
2KBvaG84RdT8PK17UpcJTOyyHN83QBMQaxoMPoHnpORpYwxPZV9v32ynDLq+zSctSbH94GgFJCfS
a/Qc8/edIIYuXUbuBp0XRaArEIiathPsDuoqNcwSFtoTDSfh2y3zCruNS+t/WDupPvPPeDTZD3qF
8hOmpDtEMd5XWMVIu1AjGeZBLhWLduv6fYiwfABwDe40FrR0JQdZQem/rxdOCCHw6+eGqAknfzB/
YjN+i7+t102FMh5xhQWU8VqcMfKdnyazBHwBkdVNEiN167e4+nFKwnbrgBB+HqtyHxFUDq43Y9Xw
gVhV/0BeUgUYZ4/yDREJVtne29OEFj/EjpI5a/tnpxXkkY0gzPkzosRm0f4F3e14GgvWc5xsKDqm
8/hhUJDF+yA5FY5qHT3HdxqULnw4zFvoXSkBvn5kYI3AaefDg8OVgsHM6QwYLNr4aw1wmLh97GJo
bdsubUwOZFX3gwKfFopqWhIW+9GXMB8k2YmxqOAwk1LRcJTXOLD2BJXCnVaVs9tiRfakKlHtycBd
JhU4BAHT8puiix+SZPVMqgf/WYGVaY4cy/sw2fDj6VIDFTM/RJ1GXJz1Gas+91xYS5HOnJB8aZOZ
8MDgwCs+h/Y22HMk5813vJNBiU/3geMcEtfnJWSL6zSWAO8WZiIE1FSW55aRjG0/NPNJntsrkfNq
yBQzhDjc5ofXX0VuZKvFZTPY1pE8E6RcBdrRWSoAbef/8M3clVnzdKrQYHZ1ZProu11CTTiP6hVc
rbhDvmJIqSNfZqn4qjRBYUvIBplK6Uv4VMAhomYymdnFGNZBCUKh+R0L/c6jp+jSne515ix5EDnZ
ZYfH/BqebQz3SmMVN4rwV6zjMjgZW/XXchQL9FXYPOTBshBlN3kWdjaO9DT96Oe2GySiKyP/OVcf
b507eMTAFTXvicyUVc545I/nP98EblMYTxTLT214ZRY7jwi9h1Lcf5nkBEkDEHCFRNqwWS0Wf2PC
XWR7+s1nmGakDSQIZGD5b6PoXsUYbLa2pm4a644mWoGNcP9qagTkggiypB7NKDkgMUvpwaPdXS48
F5qRtJljXIvLuNf+phcPlZXXSag1mnCdN/BmYrEUZe061Pt/0g7N0eVAuJb4TPopZRqCxT/2jSpv
MVQHptkQMry0mqYsLdeeT/c4TEBC1qT1vf3QK26uCneiOGkh09LPpS09ee9Lj12tD5Ljbh/s0hcL
KPmbBdifi1opcgL6i3AEEwsQxf7FJ6C+ZkH032XpjOmeJbk4Si9NTvZaHYmZntyiDADm42/Edo6R
55IcXjmGAWNfYNvlSwfRbSzIDv+ZxZdvnPnGGTPEBJS4lTlRrZuBE0k3MQ5DU0LExNK+XWxJnELL
PREPaAkWqyV2V7TpjY103pwI3p3f6WdB1pW9NuGv+1sVDWVJdeKLe5+Wdx/LQQZzzL27/L6R2IFN
m3iRj1ycs7cmgqfNZvTXyaTEXLVfQiAOshUijicKgmk1NwWLrEiH7/Rmv/a7CWSWGY7dO+EqdTn4
oL5O0+XNxSSyf6viOyuloMFeWb0idc7aVLcfDODeVnRDzuClhMn63/g5Bh4RdNnIkGPvjqHc2uNK
QDLq5Ym4DF3GzPgET3WuPoVJyW7YdcMReH+gh9FNDQ0aQ1jrEfG4/QQyUleTNSHOYzrJU9vP0TFO
fOjcirH8QptyYuyOVq3mK5pRw4Wwyl7APn65OM1X2Ll18/074j42K9pNNumL0iYZrUBpwk3Lesth
3mahZdIizzZeGFFO8Th49ZFhWIFp/O+v2Gjylgj5Sniqa2hFKXW+n9yCIoVh55N0oDmE2wdfwsjk
QJcvGfsYAjCjOSmhIrt3ajDR/GlkfNK2ePqCJkU/N6folzo2hQcwqKilefdOsfp1TLOoAa7QK8UV
YAF583PwPEJvvxaAApA3z9YBL7s5GErX5wogJuMsD1mXwGdekf5Te5VP5OuW45ntlMPFYshHsvrM
hRjtrPNitDwy64RXfw1XlGUf2uccAzkJ3L60osd4pF4AJWpcyoZqdboAxRoctA7aQW91yaa21IIJ
efC3MBVRbq2z94WO2KJtYw4/PSIOfxMCT2/hBUWN1r6ysIY0LSn9QAOCR5hqvv2qPJxUCGrsOxiR
Qwf0tKIXQZ5egUd5arDOXOe0pqCEbrin7ktriJZgcMtxPI4as8LGQoYWC5hawtBrdN99VY6V1cv2
mtG1ItdZ9FiNNEgwiOORzqcCmMlJNtIvCR5eTPGXXSWwItqfnqm5sV52H9yrXe0LQd+NRkiuCL3+
a3aKXI1M9LDahoOi7w1rorG/lBwubN5l6+C1OPJwRUtJhb20Cn50HJrgjr9jrbIqbua3/hkxxizO
EIb9Kz6YtRK4wSBW9cpqORLUfuGbVvZ0Z2AQW1sFlxt6p9MtlFymQEeMFMHZw5SD4eomxkUQFUNs
ficJV40I5hdY7frzKA1q7x4NACQFvwmVbtDGCSS1kUEAxoMcqkJMOJZz4CjzZQxLtguMPrH/umUf
s4OVW/BvzRiJZ6at8JJoQOKWPfk3zcOZkiSDeIXYl/YXnkRmsnD+4wAGcaT7xJjXugsNNb441xaZ
F0oGnTCXUkIrC5rwoPBbRW1UyX9jnpoXHDPG+l4Bw5Lo0r2vDT5GZJ7qoN1CHjlvSB+HpoQLlMen
XdTnruntGE4k0AoFe4Pt+28EJC0b1tKj3eOSRd4yIxvYtYwmTawXxIin1Bcip8ad6LDwkTurcfDa
umxvQu1tWjC0pHxaSBanbqdGi9ihUi2rgTWEIFBQIPMsaukDj7hB1ZFDqerywkEqYI7NPDzpSfMm
onMq23/mi4r43HR+b/EZf/O8sYKy2QJI4ZQLCZPWshUaCSqHoa04/bHZnIkLg6vQU8arSgtCB33l
r3Wbj2r86l6XLMw2FOfO+rz3lkIxtqI2zz0GhpvTknAhx0OIqdmRickjBjizZQ/NJLWrGSJ0NnCP
YgY7N4jpru8C1mtvq4O6xPFp74Ph6rwPqgDQ3ps80F4rqW7dngoIIfUJS7imoc4T7w/yuPECLWLO
0TeSS6aXosr/At5F0y/GGhIHIeL0yanCvSuEYIbySBkn00zc5unGnGymfHvJ8gp9G6Tv/bCSH24q
lthKRfDPtO7ZzNdIACCG9D8Am9YXBoDROW3tjYTgyVKlGpIBhTx7NTWW8r2SAp8O4r0BmawvYc3b
HFlSYQNHzLSbqy5qS1GP9+oO62Gmn8VDwC2fQHKhdcNgsLa/EewuC65ETPKBKTNK2L7Nxq0CHidY
CPd8ctLw9Lm9NKQf9hLHF671jUAXLmPNYACDLSjfU+6rQdcQeh1yvP6a9LRvxTH90c7HL/MrimaZ
qpnNcKVnKm6Juzyk0Fg0WalXvq/dADjnf0VzMQLlofLLPJ4OplBXiW7O80NLpMHmxrYvUejLvIVm
398HLThP43l8lSk4S4mfgkUkeDWvUg6R+w+2mvexz7+CxCxdtTV582uO2RdQ3TGTZiddirAHGLBb
CnrVpitJrQsVvpocGtLCp3rHIzkGqlVub+wrTPnWOfvYwpU6iJeH0S7kxvLzrQ3/c27ycLz6ve8R
OgZkMnSqspSpBZr+2LUE4IBE8RxTyUt+dU0ROWvZe4xJMrjtZ32rBmBkVtwG7RmlBcCqZhi2aktg
5d7H5x6OdwCOYZfmZaoRnHJlNC0UZg6gTQHjGon3EN1mV22OeEBQpDWhdy3Ty/CoiMZ2Iu5FvxvK
+u/ULpZhX463tFsM/+oKzOLx2kYjnyEShmv/W+H4Cezvwu1s+Gl9DMLLIJ1lr9yXWHm0EVEBitEa
oA7fwGhhJjFhfsaT4Hnwje53h0nms19/nkikTJeB5ln/UyBNvOSULOPvBtFBS3Z0Dv5QSLSFGH4f
Gtc1B4JYXecnm5SCSAZQGWiCYTc4ci9sed0u2EMjDKlcZ6v6iHRHHTh33HvjmPt2c7pbE6MGuMc4
ZxCoqj3Nb6JDm5twTWzjFWCwRNkqA+E3CsNvSsFUJdGm8WQ95X6H36xZvLvoAe7P/RBPs1gXJppO
deEkDtbSHQYKcst2oal3TygA2azykd7FUjHzpMBtXIcIqTbFKSfB/IBe9DtgxsaYnwacVOjxwJ2A
RdWDMO+qJE8WytDxtkubyy4lFfjloFHadDm3m0akHJnDTBwi6COGGKpn91uptwY8gN599FRYzlLm
QSod3BPffTgFVUIVDlse0SGjgY3LWqTH6bs2HJynZ/rkwGbZ6NZqGdPVJYC0RctgKWydLaJPtMaE
NDpbAjR3WTnUqdASIHcgps9Lx5KFzJZCx+YCKfHYO8oROdYe1CyZgajZfMWRvVzq6bhjC+7vJt2+
aMgqmeWaqminzuHdj8IKju31BzFBk2VcSKg4FoblfOCpmDq+KMFbbrRcDnampkiqt7clNurEF4wX
gjT5sgReQO/eU/d91hiHDYZoTEHgtZOIKJGp7C2Ttn+yNVx0vaXQ33seo879a4aXSIt+hiVkaFL/
k+388ZzCA+U0gDmNx6U20Bn4kywgIVCCQSHZBzIx6gcvus7zVsO18JsCZHIVx5AUNEu71N+Kyuxp
TmlCBdgGj/lHT7pKvROM+kXAX1wgrTm8VN5zcGBa6UzNlNBt7HCKhQNcbpD1MsKo58RWvEMDCGam
Ri8KNrjDcm2TwTUMaiHK4x8+oOQQ3C5fu/WAwWKQEYQEES5LPFyXqyqh3EZaBa38xr1q/+1z66fq
2r8OOH5zyw3v3CY1NsRCdhETh80RGmoR9ZkbHooY/FfOzZPNsC6FG3a/uuhW4G+6WAsrbQRjg5sJ
koCa0p3bM12uAAyFU5cw1x6YjQ71oIvEXoUptv7Gjm2R4raQOZxGtM/W6BrdSaW+xmwnq8Xzo0s6
Dyh/48DgylCC2qnuSJGBTBWGYEM/41f7vaVb0zj4K+cHUzqwtO1wzQJe/7vd8mjny7/UnLR1jDi9
n8pqTjyz7t5yJHUJUfIaKn//eA+lXJoB/ptJj6CMnJErFdjUJC8wsElcMA7oASqu0Rkck+E7CnKJ
EZLE/iRJLeJer6cVIuBiEASUFxF0lMlVL5bXnxF4RsZUa00FYjAxj/xeTfNsMo1prlVzqHX4wDfO
/7YJk6lG5pIPJuh3RI/Iz1Jdik3vymS7SUjvs4dfCm5Z2gnI+CnduF9oiasTCEXCg+QQL1nGgXrO
waFUyjxt7EoIMIqFrg3NM11qGmCkrvgCGv2sBGZoOZsZmr29xci5OViP4HJcs5w+uBaFhb7BXEBo
fbnyo2W5bCJPPVbE2UypENGS8JoS9hA855jbAiJV1EAXpmPci4mjjoK9ErMDQf+cIedjSGaJQFRV
++jMRl0jqsc8b4smyGJ0QdffLl4nx7FqCE4Qam6n49Dt+KfdDnbUMW78gDdu+cJoIFgGYhQAHsI1
22QEHaUM8sQwR+1kOTXFs4TwB17ScNnQVALPZF7QdOFXEa+K5WgxpbQrZFGSt3vsead6gFIA/qjm
7Dek2f3PK4Yuwqcl8Kcs7FBzs0U/huEZD24ATo73MZHP+BGGiCCNM0YfbMF8TnX6MUOksZf2lidV
xNc6XMS3eslQRescZ9NCl+jAgPtdzrhn2zo+NQASRR0VaFziVDqaPzWmLzgDAs84WwfB4rElPfOA
1cHav2F3+dI+850cl2NZFufOFJ9vmOJm1GolEpci8OzC1iKUYjYdLIAA4Eepfte96n8dZ9UixxPC
sv9NKXm/marX224EZP6G7SN0Q4Nvkmc+Je+kjwjwtbrpuhumzEtK7ADWaupma/RdQ/2RXf5B8mUQ
N6qs+PQT6K5IF7fuuM8NwjpM81Fyk34f3kee0Aeu0y+YYEELlHWbRjPmW7E8px5m8nusGvvm9Giu
BGaaJjji9T50mLMWkejRgCQQP4DEKS5ZL0mTan8q35IR/CL/UQaMCnPQiG6NA0/x1AbDuhpdl5jH
qd0mFh3HJhzrS00GdjEfBMeDGiAXbLeiP8RRc6p/Jci5VZSrODzw6gY1H1pfqrs9bfapw+i7sumt
goyWIwtFcIf2IF6ch/8L2W/ec9b74aBeU5W5R1n1Hnbrv+NU2ptAOpP97L0x8I0Z8JVvhI/D3YXU
GKPKUpEucaM3wtEM
`pragma protect end_protected
