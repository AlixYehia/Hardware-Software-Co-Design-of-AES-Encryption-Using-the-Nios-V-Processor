// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tfQIjOUfMLlrZWU8IMBORMM32BD7MZ8yuORUT6VQfbGkBLBZOjqFrTJdOqcYs+P34OEiF99/XZJ5
Lx9b5qKnDy4hUDiVptMPAo8oZHQq0Tz2Fe6+VRP8jLQoM3pdZTqq8yvv/KbxAzhlVzJ+1RssHVvv
OAZkvy26/Nn876/pTJCGeqxxACoHBBc+TXUP9/NGpMaebKNV8mWKE2mcRV91Q2yf6nkU7Smg5L2Z
HmSByZEvtnN4RfyEP0zXiyC6eDxubHVGiwY9PnbxDbuM2UQ0CttcfRk/7lJRHr8LGiQ02pMtk3rY
jbHDkeup/I4h9kICoYcidulkC7uP8DhIpRcQog==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9440)
nuYsheetElnZ/I0rn0n3Al6dFUP+xEVwdxcZYhBqS2fXEmYyOc6RDMtGQbnQPsqGy6CdiKCTXsKY
ZBKxJQsbNXhN5zq5NzFnJ5UF4uCJ5SsTHvI9XYlzm19Trg1TBe/YYCl8ElMaiS0bXtQbZYAGxJs2
hzjGJrPfYe7IBie5s0SDSOCq24mrOKEuhRl1bScQClOpDJX7dRjC5wVHkVS7IFwF1gilDoAXq2e3
XJtY6gySLtk2ysRm8Y+H5Itp3rk7Ff87VegcImrJpdMbjTI/M0WB7T7EO+Rz8nPZfTMvd8mnBenF
4zcP3lwi3Srxg7sEf80zaqsndUzXk1qd4oaOIl59Pb3Fz91s1ikndh51MBFr6pnHuku7B49KwCM+
ctbxfNptoq4cVJZta4qniqpuKQwFRmgP1R1WOBgkh8DQQrjTBxEknbBH0ZWgPBHF9uG3bcTX0Ojq
sAo0KT7x4/eAC23iPWwLFXDuIhy91wh4x8N5yl3WojguwDocnzKO48E84vrTWv0uoT84xGPb1EQd
De1J9DhYSepNLNUlBpNERIRhvuidy1d6t1Tzra5opBYNTR/9GbQtBnqTvw0nrIpuoEO2fRXWyhoj
+dEJhWOUjzooYR0KxMs0Z3jClACTnQnxyhQEgUEGb9LwJUabBNwQhi0NjgamJMqCsVww0zuDniXC
iPwhTcfhL3XCxwaFDiJ/WD/mUpybqgQgao9owLckKN+WmIKhjrgOeLTFuq8eLdGTEhTgfr/dF9jM
Uod0hazveaZIAKmOx4/1sHOxX6c4d9tw+A2iILQ3ZdukcvETv+E8PgDOXPNn22t4P/XXf8Xj8NYD
qUKnjrd9cmLY5Gc7r/pfcKWjSUv88kr8PeFaqDkJXT2BXOmzHVH2MRhzuJGbrtGh+QVWeI6fbI/g
NC5szp/ZTzAj15MzYnhD/oV29C5KFpssl4e5DvUpTatihDf5XzFmVf2iLjeSgPbAsKR+i8MnXrpq
KykTb99uGWksTBIj/AeXUM8TAzuoELjbGOC2gCsOnUNgg8/2sKLANPk7cFYk3GU4ynNdJZ/j87UG
qdhVGyMmLZYjt0C9h0HR3Ik2tY0iVAjtEY08SEjZTRM0ne9bp499uhsXGp7pc3NaednbPqWylQl6
561pcjPbr6zq8ku0ujCXq+XUTsDb2fTRQwPHYQr0Cibp+3EOLCC8deqiQl1yoy7/cTBN4p2jqYvc
3L+Fa5z7m78j9A1AhXMrI53DPZN03Y4TfvuYFDTlDg/9gNq27DeZqJgWoVTPzzHOY0zD+R/rWPM1
v4gS3Fn/IKdt9Yo9vPubfRWNwWkI0TL3HrtIMdBq8pWZphVgkO1pjVrQKYKPMeVa7w3x73rHIKJG
38FSMRTQCBuqXhA3qTAqUkDAggPQYRf9QVcwVvfaJkuwJsPZR6OyxGv2LFpr9xhA/LnzaaR4HB/z
1gH5yN9nG3Y1KvlhEIuNha/Zf0orHr8uGqq7xb75uk7ydNoUMr7so+1NpWzRm9V7s+w+LMw9ruW3
4JNaDnj0O74s7PEzwRH+wwWoZ8jDcNIiwRi37wXUxSuPubX/ZJiej87tOtEtITI6zKVaUSW5/MYq
m5JPIatgrL4Ov3N/YVutuJJ8DDoCdpCoOPEBGgHCRP9R0iAmeyZw/682PCGo7HrjRcTT3LG9ypCR
xIGl0jCxBcqP0tNbTWH+wBtJVeX784EDacaOSwN2KzfGOOpJ7OMJTTpvTuyjT/aVNoaf4E1GBxvc
Gwwe3X7sPnifK1Y7ELAxwZSm8ycyJ5W+wmz4GfCgH8RiGnXXOPdSQNAeGS68dQLatiJbSJqedy8+
RjYyY19J7GPiz5U3oaunPqP32qj0SO5EGlB/2aJHuNg/GEkLCJS7VC1JcCKIUuPYUzQOz2pZ4uW6
Y6qFa62/ldQIio25Z3+1Ly/g8lYX2nIfWHPpF3LLM/h/5ew3K6v2NoBmNNv6hD5qr92H6TeGPf04
DJQ2tu0582W9qqC0A6ZoY1rscqppqPwTsnmQhsU+GXf/WfmtRQaU8bkwBcAgMjWOORPR4sUQ4Ycd
eoKwznkPzsvhhPnzxbdF6ZR70R6kRR0PFIySOuL6f08beFb5ekZ/uIX/vw01mWI7/xlbDP/3Xqn8
lH4H0AxnO8X9D0oOktlbJ3FqzZgaAGXPhASpqG4BldybtRY75kQLWkSKqCCMfjVsKENdWwf5RjEt
P5UJbNsF2vaW2qdH6ohomzTg71pzXDfkYCD7itDSnLeLE4fCcXcDF30lxvLLn0Qbw826P48ToyB2
AEMmFmyEqd9S1lMKWzYTbz1+FqTsu0gR5aU4RPXZXs9pLaBmBI413wYolmIqDlJeRGGS2z8Y1F4o
vgwd7l0I82VRLR/HWWtx7TDI/X/eUmG1sWH3BKg3uwtA5JaS1rY4ORc7Lj00Uko6+1wVzKRLBdxt
JE830pvyRHvbFEiCQ6NjRt1mqbKmynfrrS2+rMbGAKV7neeaEIN5bszMLqBMinE0YKo2Lf+lE9zc
Jexffe2RF42rPo94F1S6jgbepZbI+PyDY3+90qiHiCONIdw+pSIXZNfGctdxwk0K30L4TkII98E4
qnh3MgzZEjNJgDcAiwHOoEAyFJNxKIYogMya7EtX0tzNzsqUqITCt+Y+amxPjsmF2AP4crbP6O5z
NtTklZXpW+fYfFe0JgLZzZJtzOH8SOqGvDCSCXVVaY/BY/eAHnNftq09ur01IvcjVlWE3cKaadyt
AK1lNiKqkrMKJ5EC9xur8hjMhF/tVIoOXIs4jWA+Pf9fXVpUvzslH+8ZJQ/HOUGS57tAd+Ln1vtj
WTIT6XMTK787XYoGPsGx71G+ADUVN+1F/nYkNyptOKcTnekCm897Ov3Ig52qMvB8nQT6TxzVs6Fb
jDv0nYauASvCF81Rx0fJNB2V5/4qlHAebkrS3+jEXQYTI9Z1dAt5s6ojGclpq4dUnqiz+uc40pLK
nCfWREa3qC5LvOoC1fuaTrTLSdPwImX8+/XlduMs9QannWIRjiNAZRDZFyZl742MpEsVTWe6T5RX
v019McyfkNXDjIMVWOGUR0VWjetAq5CUii+T9EcooQIufiFDVa5haCpriVmGV38733XEcz+OwNrl
v/E2n3JWZ9u/mNuFqvXpOcJu6X6sHfhvGOplyZCKnwYcLPLAwisOUStnaTs4rt0Zzn586Rh7PZs6
sRUzPKhyzueSGuu2nqm+kA3CvDbPJjWmIbRdeIPnsCodqjhgrPXbD1SKlKmLVjTrvVnSi1hcfVMF
GrSJrnZCHwGKSy/ewKOsFaKdMEv/nOks088h39Aync7UDLyyVDNjtnBWTIYmA3PEJLy/3wMcn7BM
5D8ZcwUVDsJ60hRY8FwvUoAh9IWMUvayCU2x1KDy0LThm3RlAaUcz/o+kghYmOR7UdXP9iCBxuET
N2USpTlwN3h85l5w+Wbs3+fSkJ9eqseQW9I0rl8+RLM6yw/h39WfIW9vd4uFKphrPf/Y3QguYDxb
CTxIRL+q6hhDB/dCJU7U87bzKhgfMaI/F2PrLpiPf2FRj/PK69wsXcbOG6rDSR/VQ0FGwDuOxLk3
rREYkfgkJzL6EMAViGoq8laK6V9UZV9Ey35hnug0ceUDURb8TNiER65i653ybGfJc/jualeCHLRd
fX22h+1pi+KM3N7VB5rxzTOeBJn9mt365GwvSZcgRXsHk9t/2LU0bfo0N9nAOYlIh7yht8tGlPzY
f4Xtr5HX5tnuFG+Dcmj0sZcDAMmaTd+gukxGu/6XVyKo1cyo01207oWf9IhTsPvlAV278jZ1Rfxt
3/tB1NjbMCjTQe8J7SZq5fdea5bOb4I8wIZX+mYRBVJeoebIh32r+aT0n3t4Hf1I1/NbshI3Iuga
CSSJCwLeCgREQew5z1JL/qUlhRN03YA1iTNc0EiKrkMmBLj1t3oq+FZXqd835W8+iB9DHIviSRO9
QLPXWOXMiesgSpUAyXwfBBf2Djtb0+qIH0+ux8cGS/n9jmUYBZ3kHvNXGU2Zy4XQQ1x9X7SJ5PWA
6bYg/WmyGHvqYeIF9ErAyfhUSYPmhcR99sJC5u/CDVbA5MjfFUOa8aukus/WIs31uYddJuCXegXG
n3u+vkTbbs/wmz9bc3FeIV1QDKviIWWU89o8F54f64XGjvKplB325sCgiTFE0ditvSDnopHHmLa1
72UV+m+Or9dhBKLQ3cxLFUvs2ZupIYu+2MLL0buO5Ckq7JaPhA8rY99BZ1B8C/4XmtTCikdccz1X
sOEyaWrB/hqzeoORXGpJBzwWXoZQ0PBRoinqtVaQeGz9vxLzJ98qeOsbONw1YklgSeKvr+329NFf
umqN/t2cr3RIpyNtvU0oyAq0dn7mf/K0pHVuZEr9qvdvRSyNR7H0P//fgut5v7a5CbD+TZ9HASru
SH5sX+zJArGsEu8Q5ZcamU/LEvXadW0o1oglaTHZ6Rqy568Iz1bTkSa4g5OJNB/zqKSGPgpS4fL3
adqCZOPQpnEtxYCe01JIYK5WA00uR5mxVeZMTT/nCfSAR+cOuFD1O6eISeNjboOBabLVRHTtNMIH
J9fdIMojAiPy0vxjTpuv0KdwIbLvy/mUEwNAcRQDeq8cOrcN2o6nfkDhmXgXGzbEraukQKiX7Skm
aC5Vo/c4G4kQHU+ELNGrhEKqXqp11ufwvJ1KU0XPjzPpJeCj+i+d46JiE8U7PCfKZ+nXh2tHepa5
hKcfCwpQ/+QnDQF2fl+agfTdBgfnKY1R/W4B8Z0QifNSbkXilYIYtaSYvpd+vGMosx1oEWU5vlhx
FWZC0N543j/gHbouroYcZykk5pey5zn5p3zp1/rkBYFENYqT3jsM+CCWkEuMv+qJzXoyisaVRCvD
wVE8HfIxPfi3vkPbt3l1gnDdegDJWvPgXuYAveRQBmWEIVb9k4sVwWKs6s7ma0EvdVxqdksQXCRc
chyYQ8lbd1RAS+/FoxKpVCEhfC/t9VTrbFrLrCgUHbNS7QeVj22qWqlSSqjJFMZLLm7QXEtHRy5X
Zl/Qsk/usKXKkiVMGkfc415/Swbl0aPcUDBuFC4qZeEmh6aKKluF3rL8zmwCiit04Pehwz2P6cSD
L0wH1c7pcgUmn9asVUt7hIwabxvYivFLqJWoOlZjElQeL1/dHEnz29gRHnc/3VVcplcTSRZED9rj
hn9b2iwNhoN9DruHaTEdic+lqfC+WKBWN5j2A7JhiDf5wvKPY/ogd647h3VeyuLarqK5jB6qP8Cx
IiBQoRVT1QJ5O+4NEa2ipZYcTSxplzMuEesNwne6XlYV3rnYui79apnYZi7dCRjQ62mE1W0IVEcf
Q2ERdl8a73HgYdK5fP8+4THrf+SSyIdCBwItDht4A7jemJGYkJmyF7ZZ6+zCiGJ2dICaJlH9yRMB
DHlrMRU8zKQxleiGZzetVL5Cix3A/V/15pLqR201vH6MXe6f2QdcH6F05Zq6TuHs8sJ/hPJpoLL3
tbW+zix7AvXn0u306cG/5fTXUJ1CLmQRYh1iitQCHofle8Gr8nSuglYVE2yzNAunYTiDMhuc7bXF
o25Bpxk4bi5hwXDu6VNDeU9KeyLpD8fKeflioO96avOXq7gDaeP3JsxlrxrzDI0SLB0M/LoBskkg
zJKh2lOU7ESNjgCKLVW2lGm0drXfgbsanshlPa9i4xMdLLoceuZVEpkPNsT2FEO9EdIPP+yR0ghF
A7WKhnh8o+HgMOIB+115Xg4KE4YnnrDsl1GkgZ4w5RsRB3wsK3sBGNduFW0GRNKL9LpIAKbkZ9/z
RO5ghDpTJ6tgS5EVaDmk0dj/h5rb+0i3yvjAFYBa36A+eSmquJqRouaBQ5+dBOhHsGwC5XrowsAZ
IgO5/Nbd6duHhxqu88rv/YTD8h+Ihsk7HlcGC28YlgJ2JFkGTDMedC0g82t/UYRmShP5hkWn4bmR
p4fxCqJ0Aj73gFxyz6Z7b2T66EVBlFxb+hvDe9oRUmmQlXUgeJ3/csjP4qTybGU4UB83wCyjDHsu
noUQob8S6yUSuKUxsfaqAHCudyDPjRhKEOl9RVM4G56RXIxcGaRFFTDooHOz5Qt2eyVKrG1SHwCw
9/J/FCRJSgRE3WAm9NUsR1DVTbRPlPMZtDKhUKYYqYlrv/OUw5gP9T9v179TRkLgto+7pzPOBxDx
wDxNvrLjs321CtQdN4RF+fAJDewl0jq7KP7HzvgcMbS162gSjaB1C8arDpimL2/ASr8BCvMwmih/
Zvt9JuHuUrsF1J2sEtw9y+BWCRpDSAx0/au6tr3cGyj102czzAKTvDsj/EHS8JBCcodaf/pFW6sS
fSInYv1k5Qim2m2kW6KYuYpcnNoWXaL8DirVWIB5twM5My1kNyFNG3j2HiB2LpXYZWYcih31OpnI
WQsc3fce/+eZ++i93rV91ZRhSnQlAQt1LNRva3c9ZaDorRsjJ5fP+9ksf4yvWCI/HmjgEhdpLXBJ
K7zvsmIQIFRYu80dSHPqTDHJ5ihV1hy7c2u5AkTXMqdKt+W7UZbnBTmFvkpudQyR0fVM9YVSy1Y/
sIKxyKeIg3AhHlBb6T836lG/7AF4I5WAw8lAZ+3e+gy6u2WfCLgv7H7AF+rsQd8oaUwSouJFgMrL
23k8Vp8/8y9quTTrIfenaex7TaAxPvBD9otDA9SeG+jkBb33eVxOuM2XEuhiKYw3rZO+tMDu2KBT
tjxNOVfgjfUHx8zQM5ZtnElGzGTiFCdx64rrv7uvaQXpA3XZY52WO6TEs44XDcyFvvgFNIEn3Roy
wOIuOzJM4dTDXlnHEVberqC+sT2gZwia4W7yFEbc8cayLBdBRKmn7LEkjBHru5rU2ZiQ/S0lvYxc
Q7f9OTw8vMZA46EWXwnW/FXudMZSyi36FIWk1cA+Gy/A0/PkDvCYW4FEXGZquJGWTPXppmak5fFV
FJvJhlfdnb4CsLWRY0tQQ290Z/VhFT+zDkFLLhY9sqk1zY2I7ZUPM1SFrKWu73Q7wndBaBUV584J
TfMYNY9hxf14aF1tUagyDU8VLaT6fcmKd0gzQwOQlXDvPRfE3H9af8ZNR5TPdSP9YJG0vBn/zvk0
QJ1u2DP7UQJZmOjw26WrUuBeah8yTiIR0whySq62yU4Ae5UZ6DjxG3Y/lrBntBfL7ERm/SgajU1v
AY2he4TpHUpTY41J5CPrspH95IV3XPrkv9KstUWcn1OopJcK/bUj/jkQxVIfJxtp0ie/P8qvHsDr
7e2z6fw3ZDA/tykrL23M9tfPBJogCXUVH+3widmBMlBS8BlCzsNCinPJqejhF+ZSWP3aIFauiEHp
9iF3c//SOyjxMIObav2oQ0x81X/xKER79tR7mg39PJbH3Jz5nxWOTbCcDTLLMXEb5wDKkKtQPtHb
/Ue3Y/Th6N7GPe07eheESFg2kqNeZoImKnlMZQ4T5SyYqWl4cY++3FEeGI5pcLl3f53yHZnL6chW
z7lBFvoH/Z4JYvUtj7RBEsYpNZKbrw+mhVuVDY6YvtK3zf6N1wfuIfg+f6huFM5pQg35bSaght30
d+Yz8l413G31P65ja0GtBiUExGJDCeOwNnmL+0xlJvUZ7tH1Td1UTbjk8z65i6Y+CD6IkCoEogKw
aOgiqUdUchE/OtJXs1wdyZwG6RaUGRJj6iA+VfHXT5HXskByHH+pgdeZTGwcf/O38CR46ePA9c0V
UOmKEvCQj+spDATgHE0Jx/ErnYPHienJeoOojhoNBv7oWUs0uyQ2VFV4jHzgIzmBywFEtF7h967T
3wlvzKUtVCZ2lEH0ymOyYpXt4Oy/F+r3qrLk8LXDqA2AmfaQXwmOQ+5X+//H/4vmIAgDJ0qp8OzS
RKS9+aS7rowKHEwdTvfAkH2Ti6mvm8lOXxcUsWNby8K0+Y7fkzHqjnfw9kGyHipMYXkggPlOuuJ8
pYvlzFu+kMcz6xE0SRBIrZVpL5oErdpthA0XfdwD1acrEniiNP/hTDGRt1POjA0vbcvofVpGzv4D
Y+1LhPsStJBFk0vx+jk2ANRSc+sS6TANv49mbPkxbLmJc+4S8u3p84gKko3RIFDSO7CUYu7JBbLY
pS9qK0YvfFl7FG5gbkWKjfRdrynEopz/2j2ywjC21k/7N3F7zfLR5LAqcxMCCWfLgrio4tk9LxOc
VREK7ilNWs8HjK106e9G5B18Zlht5UDviPYJ9wNVqbJdsMEDViuSkoRxD4/c+DBG1XXs91GQuD5S
sQlgqMOKQGWPKnUJfiKFQe8JphM06ftYKOOcfYXie6XlKQZGhu+vppLGQU3lLLGFSqKv/GfZNPBh
3ivZS8PiMIXZPPhGZNOhLTXc2NXqj77fxJ12ySlXgDGakondaLDbWv3cDbwSNgCTFc4i6MkjQxvE
iOqyGm8/9gkBR5qD2ktI3GXzzlCMLlxVhKfi90h+IM/U9tTVVAsFf10ehlx/G0j9F3eL4m/RrW3P
6OwDRi7keNT6Ku0eypQt8nZaHEheQHqBtZazlZTOTix319bkVH/UmQKTF6Ncnj02X4XhoSqcn8+w
zCgReMCYfBuPT9pKpsxJjYRRwxSxTNO5aaQP72Ybh5h1iTBY5bQQjT1ky1YKdcCP6DV7145RZUa8
nRkJxT+Gmp3MBEtEpmDiz+1GEGkK95aeQ1qzY6XKILgerONoBQsFBhgc2rCmV+UuMn+vuuQTiauo
05hH/sOCiz4FkeBHu4F/5Wtesvf+/YDOq+5mSBGaKR9TE2UF44lbqfYDjVVpMHYvvpXpWic65BV1
oNfBSr6MmQ5W3nLP3Nidea1YpVu3ADhVXp8ZeU/IFntxCpVtxoD7V3eNe1iM2zZikVg3IuUxoKFL
pzoerBxv1A1Ceyo5z0pLAidsDEYJnROqVnsN4CTWOUcSbIvn5a8sAovm7UON9+1bxJlpeqf9D/Au
9VtzNBpfXavss8L+bro+PkZKcC91P9gMsj2ukV+9WLYzob7TONeGvdoT3dwgmKahhmvBMVPr52Oy
JfYkm+M+EwYdZKmkSbz4CrItb2U5fMF6vuPyusNDHcjPtIigkqM7wAqdNznyLiJ3UgtxX7e7PdY8
3vxOkwn//mjW0vbEXAjy6LQ0/4tN4O0YrAFROhaZpuvSX7MCmrwLdez09IPO2/S2ohlcQeFT7AsD
77smmaUzFHx0zRNIfQtBCKt/KkrK183OmzPhthK2Tvls7Xj8I4ajB2xVOFmjLBJkMl44l/2Y8yWF
sBUU5l0vZ3UiNq/2F/3+SJakW6GcofCER/oYKbfZ+TP8uqdMgyw8gAHWJOW5roTF1yTExS5XVOvN
syRsqlIghg1QOS6MhClKRQJtePVy8WzjN8PL48MqANoV4/MbPj4M6QrPCKC0GoHAGKnJp54VE7WA
XZjfGheIzPyDHZMAzPS/MOKB4HitvRxaPkZYofEbSNnF60YhS5Zef9Tez3OoxQNUQZ+sQ9cWudNt
CdUEr3nMdLSIxvg4qmsEdB3LUvBPQJN4uCiCj+Wbu+owxQwgsEyFrG/OXPgaHJkacDeB3C/f/sZ1
TlFFuvM6pXs23UWm5vP4RVtUY9IOGbF93913FA1X7W8EicAWwCG1ZTEzOBTakpg1LzFD1cPZ5B8N
QbmDfU1FIrSjPH5cRWLWaPh/85q1+6JFkGG3T+FYDirl7PkFeU9NN+QASpVXTYwMT/knLqBWg0Xt
qK/nfDZeD38dG2sznlf52gNovKO3oRnIgpuPaImYBbdf5v/tp01NvdUbSnLGBcpfm1qG7IoYXfyU
wjYxTMI+yzBroQmjjY0l3miGhvSW1uLroctB+jjFGydwFZ14wmqfwVky4xZpEhzUJ/vX6y/90/Pc
RXc0wtFo7y0N05wuouli0RtFLriCgjc19v/qlx7j3Vr5UHMF4CXAcnsM7Eeqia+q+55XSBd/m3vf
9USwbtisxY0GhRJe1krNazWoKxISk58AgedL6B1ZD02Bx5yTqDWec7NAmf8l7AtnkNWfoZlI8kuL
RwBO7L+r5Z8B8d6NxIEI4xn3epVtEKBeeuwq0Id4Bmd9NIUVWF3On+u8vzpjyMp2ig39srfoFQ+r
rWd7bhXTtc4kryOzHa5mWMQvwFAYoNaZqgdjV7/VZrfk6TRf7fp047gOMqYJK0Wl78O10fjwa2b7
qetlAYDPQ94BMD+p7u1W8moNP1cYYUZFBWRUH0uZ4LrSqhD/gkAvYieufSXPCCzgFZwL1oW4M7bn
GAmVJnJpcyQwTqALO8CmCK2S3HPOfRE7yVoH9Sycwn9Cmn2nzDC6eY0XpcKqYKsnUcaXd6uA4OF9
bgoghirsfiyIhD8pdqnM0kH6RohfHY5CtL3J2xefu3wKK4AUPLOIs2kN6ZL9c/cRNsET7fgdIc6P
RfXSdlPtyVBDAg6f36f0KNLZrrl0yBDxcE2fgG2s3Keg+n2jnOHhdnzrV/7iqHuc1vSzO389/fIe
E7w6rIAoKk+s5rfub3e9m9wqPem1XITRvYJece2ohLy0rfHin3HQY7vRcoL7t2s119K9vWCJ2+Zq
dJEZTZd7DwcLQBlbXiFzqM0yCePE+Z3gj85sTFxCiX7aE2FCkSDhIDCSMuHOKdggGHIv+hlaeWet
/mvOtUDvuwnJ9FvjWyn78L1xprWJCXof+A7TWXgGUeyiJZiw/MYPTk9z02oxWB70AKGGUoxPfWf1
t5GXskdy6IOWdcPoKRjqkdWv6xXOyYvIL0DmbPfEdL8HFK09a/xnLDDK2wpQ5TvtosLVPg9xrRlv
P5SF58lozXSWpwBZ0pL5CfDzK/yN6dMbMpTKA91+yHTb+SzMJjXhaQO1mFQ3U6YRgG2DbscHUHsz
0ae2aQ2f0JuZpWwsvpA02Wwea7i7EpiF/vndm8ruPqiplcBVpgR/mwM3gjElNi03jDdE76hts8UG
79KeqHULQ257V5ji8Iau+P5PgqOVyFCGJMBXxtVu5bUM5ge4jJ7oDdXEPWn3RwcQttUAZCVeeAYv
C7DTnsdm6Wp1ORE8iSmfQKC0710ax2azUgAM87XHAEGlX03Ma7P/AP2t+XXJnO/nZUkbkvELYBwn
Ds2yW4zhmQCa4hxy4MZ80zlyX1htr57F3PwtuI7v5aFJIsPcrqUV85jn/lqLFreb9O4iPN4pHBFO
32eloB5+CXT3Jo2/j4UiAqrwZj6VJ56ql5NwZ5f9OMH81+fBi7lJHTISHr1x283KVI1vyuRUIpOs
/84mr46ltxPCPaJimsEIdk7PBDtzLuw4NHgpatwRCJ5g1pzJwY3uKNyoYxWOWFAhV3ReEhy1QYVR
VNeDt2C+n2k6OLg3vXusj4ER/j+4/P/WstGRPDlKqAo5eURcU1aEUximeCt5YrAVYg9ekyhrsZZK
DQElHvylKy3XcvzvKLpo5QN8BzOxGVUg7/dDMjTkM3grwxbd2I54HXdkSraV64UrREQeCBg6v4nN
Xuv9MYh7GBPZiMIbLkm/6gIxAd8vkg8bGBGxFykMbGhsRfHqdraNYCT38NLSZzMKV8e/rEZmSzCK
tg7B3KFPp0XPPep6dm/hYY3zO2XWCXiSIh5aulJyHeO1vP5Mp7EgZ6FeY/eI2rI9hkyia9JvwCHW
ZR48jNh5DL+HAT27Zw36Cx6M2fgJ8/fXTTxOEwAxM0+SkLTIsCr7FDLrSlS8BoCg4gt4EcvRtUVo
Tv1/W0HCqoKn/BadD0PsklT6GNEW1Hd1oMrCW/+tbhFQKy5cAhvPgbnTDlbtHQa9jhqzzaZPGrKU
RI6B8WasVSJbznmOHIwcmiYXEXKQsQKwfQ/M+rV7oSx+PzFQKj4lZFoDWD6sWctvPthj+BsiDRnu
lMdcSlvBtMGXkkPYnNU610pzs4Fc4hmVtL+HUR/6e8t1UzTEGPJWffRN0S+efuhk+3rtdmnLPH7Y
4Uie89tm2bsDfTPrNUSfNh0FZwooaU0AJleB1FMp0Nb18iLUSy4AQgAVwq/wbgylegEYEA7GAQwQ
bkq8/zTrJj5ELMwt5IZOXsy6f/ofGcpeOj4oveFQlX79+N26v3XEuo515nY4I0SVPV167JowDgu9
sPKmwsR2pQS/2f0jsIMbB+a+K0zRpRkJ+9DIodhqMOwn8hio4BW/4b3N3p8RXB7xw8iB/N4MI0z+
LU9YRRoAYF6Q3jIBAvlr6JBEkfuPiRDpDVU5+m74+aoj6SyLF2SLPY8NjFAOLn9jEtj3aFkqKt1O
dCaJkrhR0X95Z/WCvKoW/vyXmjov7WFY+IZEUPO/Jnx2P2+WPCOTNZbdOaLfZ3vNSVQvTgLx3svX
C6RFn2gysfOj17+RQ6GgV107fdbvZg9JnUTN3Qv1O2bGINQTlRNFrM3x5jQLpED61Tdd8Gf+0Idy
z9jtLzF5yyZf2Z2DFVaZDZolfwfUn7MURGec9nOp6i1SWXmADvSt2PIF1N/UBkNw1iCM8AcRZFF3
3PxhNv29KbA0ZsiNkDgemin+VLGi+AgTscc4MAOqaIKnzKkQI8ld3YLJqqn8+BA9CyIo0RgIcux4
h29/zUDR5nd8imKwndWtqAbdkpuKJnuvB8CAoWsLkkXVfbeSVGzd2nfsimKVRl65vmtAgD6QcYZT
59pV1Rf8TrpgRRnXlkWFgHRtJoKVVES+Qv2O7ecBRgwhXdY=
`pragma protect end_protected
