`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZFWkQVxpweyNRkKtEoXFytl0UIERwy385fGsUmKlvLxnrM5VTlG9SUwBFOPC4Tku
I35PvBOPgqVbWU8jYsb2KwMRKUv/AJJDNQ0agM/osR9E7OS9oHxu7UDM2nSXd20P
5mfEgZNZ4iq3LYYBu4LOKdD2yS13uUl6zQGUHjYrlTE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11152)
F7zumJnmEA4798oXWy6mmc44Aq9XEa6qVfLXmC0HeWZBGdY+SJA3RC38xVbhIDWV
7W9a/dxTyvjKdOaRP69qX1A4JbsU348I/tWPawq4oOvQTPsYyeGzQbnWRr6b/zxL
OImSfYin+7EQpT8XLEHO1khYMUIN9ftN3PdwvB+hWL6etrjF75ZQlhrm/ZOplP2p
4JudTn+Glz06u6FQ6C8OsMlRateRW5CZ8dOwLEieilsyIYMMRnKDo5JuaF+VHEOS
7WQjv87LuYsFPJBGRntoy9M76RVuWs+/ge/D0DAYq+wuGrtLmkh68AgLwFps0CRN
MTngx0+7EfTpCoRArF8+cMkSrHHIaa3AAZID9yfPH8hdxCtBtxKGfv+LdKLGrkB5
qHztW1JxvIOdpX3LjoGI/h2yimMec0jKiMFrWb0F7EAJVfCibTKF3Kue2X69pzLd
6j3CAJ2y4cN2wbRxugi2NnHO/EOYATvutVzEVJ5K3psYbrEmocgn/SzjC+X/VPF3
8HiYwc6aBKFJ21Jt8BoDm2XBNbKCYN3lL2mCNA6tZMhjO7NmD0BK68WkEYk5/i/v
1UxJcegtD4BNlfFeAeJueg5d4hvEqECi32kfAxWYMxBWxS3p1d9JY/+FubBhTVex
DtxjCGm4A/gAYhzR9n/wTe7CNYyX+AdC9ISSWDLj/9sBnDpVU5D3A+cyjPHDM7Eo
JprRz9cBNNuAp3Q0kSmYc3Jy2V6+ibIk8XncV/eVkeXIFhzib3cb3bKNaCKaDSGh
5lRRFbzFFEkP9hVaAw1nFiR00edYJs4R8w7McDm5AHg4xaozHGsHOoeDjuWc30i2
0NqN7Dj+xISbvNq42MQ581W2cEXUNt4/MFY2c+EFi3G2cT9gFfleDTmAv97cGEIJ
Jqk5wITBq7gJer4l5un7u3ay7GjyblR+JI6C4HQVNscS74Cgi7mvXRWATkGm1swy
/yLwg2DXrjHH4a1LDETGLtZLE6WwPWOoPI49Pf6p2x4l/JXh272sQKzAGmEUzoAQ
bPg4YDC44UtFx3eGFZQCBYxuMdVPF8DaVDoW4bIxbrTnxf96c1Yij9QNdkImT1UE
Iej32VtbGnN7s9uy4zOP482o6aJ/U7gyKRYDK/tlZHaEvnvSq8KNGE8NcrY9RRaj
2ykaqmnnZaZCfjuVov/hpL6FVv2ITvk2BeBg6Z9oCouZwh73WF6sK2CnV4h5pb4U
QoFKzV49Q2EODF+VruY1UmhQY8tYlS7m1ktJAQRI+glfZ/TBXAnnNtorkolKFaF3
lthsJp3c6RaVTDRtKDlBwI4PVjsog1r0fZi86j1HsZs0ob66/YNLreepjopOUQOH
aNbTy2naNoUfDZlq3/18eRSqfulM+spyXYAo7AxidCJvMrfrafgnygm2DAhEID0A
U8Txpb9py8o4/yF9LzyHWhf83Ioh9jhfceYwZlXFkUw3Pwb2iv3WkzYGobWbiRw4
paKsviQT8C87whYiUbH0W0tUl340X6NuXJByfv+jucnSStXTfmP64QbA4WSPm611
z+/cFeOW69TYsI2JILdf/Em8YIgK0ot2O0nNDIDAL6OO3xUxjg9zJ4rJoem2u27w
+B2IVeJcUzhYWCWau2bhj34aZ+FFI0hFFFvhPen+lDBNh0QUQKoeq6OtzU4taosz
musGHOGJ3EyPE9dVqmaYXHHiab4lIujADWrRRsbM1jtYSjCHp3ijgBcbJ8doQgqs
XxDqsoiTwgUZOnE765qoGVqCBJNQcaeU2XpbwPy1CfgCcWx4jCWB2J1agX82pT17
XINzOMiOKuzFDUIv8UGchHRqS1AGVF70txfwrwJ3WgH0J4INqOLl5lYwSx1sixer
Yq05VFt5dCqDJE+9mqKroOlRkTlEvEViwnqxqEXAkDcF5aHxbuaFjwYPwReQTfk7
Bj7QtiuBc9DihV/QDLjrIayhO2QwvQd4TIBeDkDlmMslt0iMJ3pOKlTAR1bhrzP8
OoLmLzoN/GeCwpK7kJu4vNUVPdq8pe9+3kOdwlbbNGlMHlB445dWkw7qcmsVU0cn
DmwfWXquAhSGMDuwscuBvnhWcp2H7RWBNwnDu9Er/cRQrvJ5lNwHzk3VYW9DUNs+
3a8apaJn0YX2eYbg8w2deyTJrna+H/m7d60HLK3VX230Co1E0TE0wUI/0B/wEAt/
3/zgfXu2CTbzkKjxrdd5QcSSfXxC1MWhKqrvh/lEFxHE5IGniS801ak0UYMN9FCa
dTPaZW9NHa7lu1p8CJzU80SrMZgDpv/g0W5L/40wHD7tOc3E0k0Fy09Jv0NibZXt
hJuglbnIiMo+eIdG0OQPliAOTDgs2ltIAkRmDEmzYvCe7PeEtH+Q2nx+DIDnHd/r
Ngm9MSeMIZd9h4oWTUVdVf2xJl52WDwGKD9au+B8eAMdu97bpe8FYbHoIIxdfqLo
7imrlb+FR+ILIZ3u3LRCw/+f9rjCTmRzMlF2d5RPjFcZCI9fgKtMRgYqRK0tOsa3
WtlhDRyYc5CJN9N7oLB/XEy5dxX0hrw9VikieX2/qJIm6hlrqSFwH1BU7pa64DRM
uh+YLcCcxexZ4cm5EdhzSGbvkhqHZg68ONC6VgnVT0JKb7Aiv7bJRgpvpkBi6C7x
sv5uvwbx8mqenO2YpO370//dJ9Dher/VXuqxOTEiexBmnYBbHTF358nnzx3H/NQ8
fLwneHhF+6CxngMpop9i7pkpVqSdIlsiYnYq/eZ+tLi4KLXEey0nnDMcPA54pzLB
Nj6WWPLwsCFB4ac6DPhsUPiQcsSZajb034HtUSrXFsTF/njng+8+dAWcNbcNnNGw
PbNfD7qxjEhQp9yuGnmCxkOoIlkUlUQyaMyZIPhZymbbcV4+AuQp7Plls0x7atE/
pOR+dABEpzY2rQvI0cky2U/50wGz3kFUBZD/O7ENzr7Bd9ULDxF87x26jYEsN+ea
t9cp1eWxcaLj40JOuO1AyK7FaaKs6zP2LfusLDAvI4dzGJE432yNpB3yDi23KxWD
xEcBp/6iwp5WaUub96K6XY5mg2VzZPOi34waKLQSt+xVbkQrGHsSPKu6MBzEcY7O
zVVNZ7Zdo1/QI7bOuAf4682za0aKBeweeKN/h+t4VT0ybFTSaqY4pnLunzYqJsUX
q0oaAg/XmLAwc6G1DlWIdj3Ex+QHlLWcMBG145yXK2wvlPWyU41zOgkHjLBBl5t1
/qQgT/KVV69pbFKYwFoFuTlH7EHBlNeLbClUhwnq1iXCyPdu8mg8FLehv2hywWp7
CaexiSut8NWVrZXoMwcPMTgCO3Zm2mN+SGGZ+QVjxwHaafGjYr7+qjrmZ2dFjKpJ
mJbrDOCasQobBMo1EiyJLAtZ1GWvnCEWpH8exVqzu1PdP4LoMDqMgYTLylRiZlOx
9e6/ry1A5YFSViQSkITAjwgOaH5nCSVWuEqoo3Nbhmfl+OL4AV2sZvjuiITxluVe
p1DVkebOjJ+J+aIwz/VoCKdfQYVI7YzoR73e6LM5jj97J2KezjcpqdMlV3/NXwTJ
KqcwyJhmL7w7YfAwLbE0yytYVzjYQlyCCxmlCZv+q3dNDECEPoFLW0VaGiqrDW6d
wfkvyAIcialM2fvrcp0FJpsM2N99nz6IEYAx112XKXrUCLpI8H1axE4yvI/e38JG
j0j4FB8agjamZM/ZJlxiJVn+7//Hl21Ddz/hE8lid8+1xsC6EEdZ9pgaLJYQbiMW
lK4tWNP0zh5t3xPh0CjrgJTbEl3PpfV5QblwCc4t6V3OvGw9fqlYvkHAK7Zl8C3O
WtKyh3fihvnOJdbl45gt+PUn2+F+0w3v5f7fHCHMu13RLxz4Y+/bpBKoF4t6WGM9
hrUGPgv3KJIFfSgi6/a95KgcI42seX7EElbbbHZcpbMzswwrOCeG2DL6GQfYT5zN
HT62s17bEszi9e7V46vlgAwtuZMInFcer/jk74RBIjQit4nVOsaBrkt1N04UThcB
SKp15lTMbn/eKJ8Tgqt9paDaNI4x058rgz2wyqEALRbJdX9lSyHznqvzBQ1UC0pM
/9EzedEutt2iHYhJpnE3kZtEDfXvyRw71x9YiQZnbnA37no2Q4T87GLfgks6LCNO
AynWohJvjA7yYTasxpyS39AuiPwpXHpW5It0Y0xcqHhB+9JznBPeGou7gYW7A+y5
719J7SNCai5g+wAfLzhSIST0lO545E3NIveh9Bj1f/MDJFOx4LtfG7RZJxrPyptU
ixUK4nGwSjapr8nb9DYDqC2T6DuIKaz2uLgazTexLU3VbiJ/5Pl9f1gI3D3br09p
dCg/i/rqmSKz/3ERUuOOqoD59Nlxn1cqSXUKQE3gAJRmHiKuvJR6enLe+n2Yn4oT
kLjz0vofvpyd3jmjsiZxgtI8G1rfZoMARKrQVbPjV7h985YHiGIWPMCzCxfMqT6N
0PtQKqmXHtqDxZw2H81F1pfoNKVRdy00AT229amGheZFjczw68F1XuYTYm4kSlJr
tdrZqJ6aMY8ESs4TJXUbKeqtVepj0LwqjOSxSFb1LxISH/QTV1d0ptmPf2jasgO/
J8wSYU9DPQdUJiN2DVITdaJQalrsR6Y1UddQXiXJCoTlnEbD1DI8tTXmYFaaqz5c
E796xkHt5Cqc8U5aqGmzC6rvBzYmM21oicgKmsxW2tVta+jHlZj5T0E1sZMXlfEn
SpmfjqbSlvve/YMOBZjlbEOXUY9V9kXql0Xa6CUz+fvfcZHWX1d3gON0i9SULH3k
N3tNkO/Fuzum5HLya1x/QkM8t6nkzfH5iRV6cNbxkQ/GKX8DueZQUT14hEWDtZjk
8Ksnhp3+tkCEyxYOGTBTu4ZjGtYXMaHbbcdXwmtu5fL0fltAzwJkSr+jzMjztXmk
+c2GyXDy/xJuZvXW/7EX2y7bdKMstcngNHk7M1H0qnVdokyVYVx16wqpFunKdqOw
X4D3ZuAyTp/f+lrpnpw3cJV+v/iu5AUM46nH65wUoUcAIYgZwazdLLq5XyhS/dCn
1k7mDCX3QGFF36PdRs72L+N5XWJB4/E6HH9NwA2bXsATczmnueOf7PChKNjMrOe9
xADQnag/LsVHNguoNK+95bOc4ukFJrWPbOY2wUMEgUrX1rJYlnQAdwWkrIOYBVFG
hnNF5gmmbUuH/Ie7I9EtkR8N2PoEuLwzCP9V+3j3BoZaXDvgrJliZ5o2jB5h2JZT
HjRLjt8znKx86WavYpo8AlUAeP0eTOqgx4AlOk6yg5plVaGOYsJwmvwLmkXIo4/8
b/Jr8uECXzUdWRBbuY7EysAoonGP4b64/uy2QXCxl642LYf5bBZo1UfXytI0J5lV
VG9gRN70GJYVIHg62ioIGc+tU9BQ8TkcT+KDi+E2OUEi1CMAR+TPUTeTmnW5e1ae
H4mGPdqMEkJM6qZ/K+13ONrgqp32ASV+mGaivIZWf0+vttXxn2lNhQ6H6i5yHBSG
Omg0UBU6pyFAzDCMM/SXkR7hoIZXG+CoFoV60Fy95XDVkkw3tFxs10nZPkHby4oa
6gXE8lGxZCm4MllCtVd13UtTuKe4x7k4UxNBDgKpGR8UZ5Zuvqq/vRzGZ86iDLYU
1EGvQlDqOQVkkMIQ1RfLdFsH+H4hypxWRoYAY8VbM5rnxC2sOEmp4NRz7cb1FvpH
F/FNRruc2W8JKEnMc3SJo0dblVmkqUTH7lh/A+a/P1maO7AAudhpt2nRLoeH4/sB
xt1Eqmr3yyoFrp+XDZMpV9zULT1ICmP0M8SaXqN6tZBQqTOgql71QQTMMW0Dkmkx
+i7Gn0xBs4UAWOewDYE6Y3Im16fx/lVpCwGO3jx0YFC2fMdY3xENpcHLnjE4idfD
6kUqAMWxww6PI51NEL8ZK0RgnVRGUbnDIs3hfqvbfUkLI++wmYlfPnn4ct5Uh1NO
h9m5+iW2YAM3bElnKugJ/1MdWskj0pQIXAup1XnJ9QGSYtjwD2eeCRcb9KbSfpTN
aFEctMJ265BNgtwLCowMYAC8zVZPpZv8nmurQRGcfyB8FphqdkWXgRw8RzWB83Ca
GSIJm7voE9Qbgt/IYzOWeSoLmxiT0aViCo9XbhqV5XAETj1nNjIpoEJi+rxQ3nis
SwDRmp55u7hig6lbOIrMLny/UVpDg4xkeVnZqrhAYt/g92PtPxl+qz+PdPr2DrmJ
Gk43BMBtypj9B9M7QdIZhKolrDtZRJteB+WwEEz67XINhhAW8/0sxCF2EwUABtWt
3J7Vle65ESZEgmAHxkyWdi87Ygz+rtkJ5XVg9XKJuahKOcIYAqBgd4eGFBrq9JuJ
jsXDxl5dfTOo+xX/vDP7u6xgOTbhoIYYTiiRXsXpwvs3gKJVchmn8U19VELVHVjY
JzmY52x4EGwRyDBZZV1SSSLPSmgo0gccPp9fp5CxyU2K0FtR5gcWJiUCTfizC7Cg
Hqz8+zW73fWa5kYLdO0Bq4dIkK0uWl+6/6zu9XHGIZyF6WkBDirB4pijs+sEjzBR
Rn0jQtCe8lu151WPqxjDXro9oF/9/opxkCzZkaADScX2TWe3y5c8nTH2y4PBFcYJ
QIgQzIabkEeHxBrMLtLRckPaAfretjB6iQm8EQ+UcfJi8au0tYT2aYwqLUmqFVhj
tOpoS/USRY/zs/cP2HyiH63YZvlRZYtwjexmaQ45VpAM3FZG1ZoPNARmy7UpRmRp
pH8p4TdBHdl2oE/v5kX4FxwVtTKNr9nAAMQkuP2vyYUdB7kANUkTH2HM1onELx0+
gAiRMU4elafHSesQfozUujlxHz4KlAdEOMAcXbr9lXDBka7xswVeXyAGFylGgNHw
CchFZrdoeB3etVBZS91WXAZq3t5fqyOwMmF+fmWZva0KrFfxllRYoo2kSOW6Zd8F
dctp0cYiC5Ci0hzi4l02Te56siGAXwHLzIBPjbIHRSjbowXPFyUcmZJuJ7TJhdUC
crzYmQJck6nMFtFdvDgqchGLl7T604YzGb/nGAwYG6hXgdufFQkvwchtIU5BkpEn
+G8oQMGCx0fIZjQ4C+S4GIAssKrqWjn/+s6n/Lri0ahj1pKEvaSfAdupkyPEuSKe
sDDpygKt+n2vZAyqYNslXNQjwaYkav8xq6fkR4vR/ZY215BcFNqzJqBfTydJw7N6
Z9X7sYY4QyrRvp3qdv5EODoSlY6DV8KRwofDJVw4kql+5sULIoFrPDpnEFLKEglT
ZuTNDMB9sxu0ElNuPEveNeYnQg7r5dXpqyQSW274q0yRgoCLmxSMLWa4wPLS4r5s
uuhlceJ2yy3cJRI4EhzBst6KY3eWTBXnnT8K33/BgiNKQjqXQN2fQRHTPEHLVrxz
J5Q9jXQYHKA+jm24h/91BLHGe2JMRyGvCS81gjFDNDSgeAMjvzwnSAQOSo1RlCYw
6ZkpiK7QP44iZDjmI85S2Y9Qrfs2S5evvkTLz/sc9rDw/+MD20fBXq6CRqC08eWR
xcPxnlb/T8plAqxgAbOSjWrQk3c3xdL0TBQ3UGYNd9hVRucRqwvkbAVn567aKMkE
myYAlAQQakoMFVzWy8WCth+K3FMIj1RqhClD0e2pgBIW6sHIrBXKUxdYiTzUdwi7
faeDVBuLdiN9nPHfEx5rgI/kHAgv5KFH9XjGbmFA3z+qs1APzsU0jQWjd5k0BsvZ
AI30gVmTZxryRV7UAsz5NdR7vVM19gyVwkEfgXVPr6nwJUM4u6Xvl7xX7fTL2tC0
lJwzEYkIs2KPA9ftxrQdeHVs+LJQ6daMMwg5+jNjEZa+E0P+8fI1YtmEK6UIgWQ5
2odTPhScFQsMeHk3hmDC53oTnCW4q/kRx/niDkhR2Pj+MOvBdJdl4gyvuVrXNulA
rBwGTTLMVESpOJ80aQkwu6vTnaCoBCfxnk3aWbecXPP3AA7r0hdS6oDFk+frtR+r
vH7bUJ3movYKWcRiw4a5R79gdb+dOw8q/z8D2rgy3Bw61lyr/Y0XtfGL8x1+sJ25
BZzNh35NhhHfhXusgZXCqrLFHi+bh70t2OlpXR2mM5PIWVBFTZ3j6TcoSp+1w7GN
GAnvoKBl039Aad1CgYzt8TeKaGa2ZSpF1k0v8k82NOzadzlcE2bd5a2MKDd0Wpka
noDd6fjzukmyX6MwMSfx75M4aEXJSQuXDPFmzByyR4NN3u7dcgLn6SD0nn/t87d0
92cWcg0XgZQYwoY30+FXGqgOdEuCr7Jab4jmFGvXMAZzHBVc45sQUr5oLRcMllrU
MVynZ0/Q7qshwn8Mwi6v/eauYcMbzGecF8/56mCa20QFKmVf8fivJyEO2oRxq+Iv
3o2hkCy+PyqESqkiry8nGAiTwXzZR8j1Te/BphtMh4lwbeW0QKZey8vvIQ0UlfQY
jmj/fj6oEtMmFYBiDCyJIqk0xILnrAY5cbbS/PnxIuNVEjIpZQKS3iP3G7SZGJrV
hqeqC6UpDnHBKGnzIub8qmHoxc6DrsQtmp75GL0l0LMzIV8mga20ypucByGm0+gD
ls3cxSkW6SjZVGD1oFlqv4DizjTESuYp4UaoHjQGjT8aNTJvRe/8dWc5otrrA13z
Vkjr/MFAqMQd6vwYgOpA5CFxszL7iMfASYFTyTS5MOYSk5ctvSkVa0IAJQ5Og+W4
MXDOC7A5rlMgWrchuBw97sGU2tTKFbsuneBwcUt9/8hvcJ3kCneyD1MOxwmPv+ya
+GUQvUgeo9+3cv+aBhuL+4QrImmJP9+iLN68B9zle4PVqurSyUi+8oat/tbR+6p6
M0rliWuIamouZX6/Hf6sLJ7DWsxKGRK35XefXczjyZaDhau+NLbDfZjqQ7HlL3HC
9Iwm+L/K9w0SEp3SRfTZAGpCc63zwwv7RqMAXjbowL1tN5DprcoeaeVyuvk7JpXz
cmI+tu1golJwButxVVskQCrjxXpVf2rNt7FmhlfRgWkfNn/3Rzfv72ER7PtcXQ7e
ySeVC7ubBE+me6cUDpyizZywVCXI5TTGcBlKdPfYLCg1t9s0AUBG3AmJQJMypNOv
vqut+ZwspY+OFu0dYCsMybVVfvJz8USeEqs6Jeh6HrwgvtX1RWlN6JxsyfGLQz/9
luI/ulr3mBc/PxDDI87ymMzhN7Y5LCSX0fO1ptd2f3K62erq7g4jogpTBoFhfP7R
0rC9FOoaGkdsWBY1sx+O82Ufa3g1551qKk5uq9tO7g8AZa2N9AoLFzdb42AeIc6R
nTw/OxaLS4aP9iqVIJ0DKPp/h2GWnlpjxB/TlAdXLaKK3vvqpx3KSLPeVARHSPiT
zU1+xWkVwbBZzKcqtXM6RrvP5JyMimOrhR9RkiAimgHlMZj45DDDF/zXqb731emI
2aayITGsCLVeuyfCeU7OnstmQGFMTOkSV/Zz4Biqdhn5cVEo3YTs/indziLYCxMk
kBV/U5AnMy4WaBw4YDC55EJXk+cWwD+DMlncSCIQmhwAGGBT3N67YfK2VSixutQ2
g3G0ZZTObds1hdS8f72eIPkKIGzTWAoMbRUBIT2P2mKD7S4Cq6fUTu3XfmgIZkS+
TwUaLW1TFWy+w1JP+6sfipua+CXA3fAIhNWQ/20EDhEL3yUrVfXXUeF8kC2tpV/K
bqqWTzmRKOB5FzlFJJUWQTFHdnGFSEmHERXEDpTDi2w4IPpLF+CJt1N0Gi9DdjdE
RC9anFBy32jmFB8gDIVAoaivBqNGv43EQPXv14Yy3zSWox4RT/o+U+OyHdb+WfI/
d+HxKqMeRwiSWMgYfr8i2341zuJq4z8pFh1tvL61lhyl/991oq3lN7foHVbEglW8
Ob28mi9vM6OI1zTingI1nvCWJovfHAgLbH7Ec79AyCfya1XzNAWEroLkiae6Xxcc
2nyy05A0GBSP61pxDkwR0BhpWAhiAI0fiYQtARAiKHryabfJcxzh+UOtv+yD5Eoz
qkQCDTPTI/q1yThI4k6OG29W+bUMc9GSOQuCdHCuD4Xo86Tjm2AbKyv1thSMfZeG
BbjHYkEvz9uBBc1wQwcO4R7JqR+nsvflZQ9hE/PZJitslSZLMdbyy/TodcZulOgP
JEhRd05TbvGgGVHBGszdylP4b0MsE2D+tRXQ/LcByGpzMHQkXNzkItSp99GtnsM4
93UcXBzFIDQfWgZ3XlXkzjnQ+WRmaFVSY1nqKK+Vr+NwgkNDSrK72EGDvFSAruMG
+yGAys6GBwsGTJDFAJPTUUVBgEp1CIWaCT8OHajpTOTTOwxbSY8sJsrmtmT0PyNe
Z9uhRWHFsZBrgWLBHZcCaniWabpJ+meXF67ixezyM2va2eVwOVw/yESSN7nNdRgU
xtWbpLNZjrdvxAmlTpMm0+SxXQPe6AsXes1iF+Furap0DIQEc388CHkhH8Iw6PvR
tpKdzbm7dZrXPLuku3iakAyy9oPLhqWL/mB7xabveIvgUrs9e8xPQ5vnN4++4g7C
chafAaDGhrec4UDz1B5STqOFwG7589SPfR8wsTjDxfvgXxCHYnH1Zmp7MBMUoOFf
jtvivQRM5lrcNwXNR/bElvv/nQg0BLfWY0HYCRwR+q+WLGvOfUgxB8J6BO7B36a8
vMtb8oWrvtPf2oGEs/2QogrCqPcaI7cmOO81XJH6Dd/MsmpM9fM+En3Lj/V9pgwQ
at+kt5lRI+gMvp/qGYTYNrQD+H4To2I7Wg06QcZGrBPRRFFlItpmllNdvI2QpApd
ijN7B2BkYAuZX2cMV08wTjEv9Bik8CF75KR8RdYrYmIKv1434GEyeOT3DPwuqIQm
42rfg+5s829rLhyFJIGYlyGUSWxm3JWsvX0m5Gbi3Nzf8vC751f1dnO7AS3D2jY9
DIkvxj6zYD2CGpxoNDquj2RRyMVHrcdqBfWvyWcVLHZIP3kvjgQHxd9tASRJ00my
wV0CgN5MIJYPvfHnLUL1C8MTqS84sRNKK8nhODC8k0836pbUzHMnG+EdAyF9doVF
XfKfteCvVrHhdTGvzrPnpS2n0zf5l2GyuXfOITXiMPEdrrpEQgE06bDJ5pUUbdas
t8gl91ML5gA6XRwK1PE/7pAOlAyxfsqJz7LpAEUX+mIKI7xrl6QVyy1StA/LjQkF
TQArlAI7Jn2IPvvDVzjYno23sU/qTG2F1cDB7kCRFA8YyQ96bI1ocre+j4HrNQN5
rR6UO+1U/vV5YyHRLe/KEuHPKkJDMH6Jq7DKoVh+DugnzLTihsiBMyqctx7O9fNr
gcbfu5sE0w5Al/enSMuml3/lDM9N52TyT0J9wJGC2zuc18enPSwDKxDJ75NGf2Sy
Mi8Ic8tI8zj8GKAlEmwKj2t/chL5HcIk49oe5PiHzPVNnNSN6w5Sgu5ku57mXnim
+CUK5BDX2j+cbLPB0+7QHTq1MGpbXKVJn92IkwkcrUeu4uIOp2WhqT1iHR71/xdH
6sBXTMkzWi093m9Fm1h1LZiwRIt9UrbO6xIHVsI7CsVvTado20sUYMmTaOogA7rK
pomZmMW6wIv8nxYf1LXc8mkdWeUyZrOwi+FVZaE3P03JVk8dX34fUUL9ZmHpYU6k
MQghUOJhkfmSPz2F8ZGq//aQ9YS8amoacsmhyYN3mF2EfhrozXdS7QOLc/Lz+bgP
bC67gL9RcyTU4tXlfVA46UnJ08tHtyOyYQpGnvRIPB0iF3IyPAko2InZZU97eG3R
OU9ryKxKSi21P1jbXn46h3X8q4F2fN8m74medloAlA4yVTWJg1aHKJLL/rRChgGN
V4Ln+Qz1q/s3o9pkyyj8nPJzGMSsoFjVBSIgZjw7JRtQbDdD32zFAAhN5RqS+2fl
3mYoqbDRekqZcskZyo/r7Om6qYWFcxQesKMnFXLFKQGz38/r5RRb2D43r7fUpjc0
WY/9D3sd1GOuK298zkaPGFUYlL+pkgBnOeHSeQeAcpvhDI8g5O1qZgY8I6YP0C4f
QcHfuvR9IdurGe70+fe33HOzzunOkqHQZIVJUavbbl5qkiV6wYf6QRmey3Es0zk8
2MTh8TVhZjzDyuO7EE2cn6hbB+HMtz5PIHVen7Kz1tW/9eorvEiwtxPSfXT8aU2W
CX3PX0dZDpFpyDwu4tWdx9zezIp0c8lJAkXR3XmfjYx9HZLMhFFUr/Tl6G6xHlRN
RdVoj4MzOjaj+XXLi7etB+tkbTY9ERISVm+4ayNiG5icenimTzgglUcHMEfa36GI
O3JG/hHJxmMlR9+qan2jWyvQWwNXCGv0I7+aRgafn1kXZwz2NGMZvkE9XdSq+Wjt
Ca0phxvoFOKbwj+VFd35lizKgysdyI7W2ixcArnf85byRAVI7IrvSxRwx6I5sjUE
yQAtw/HMCjzFSS86aeGYgDdwFF2EdlykmNTbu0fV2I3mdJ/LWS5ZFLfKtruP2vn4
KNmgmEobMxbdcB8OlFmQSnKwmtNm1VACY2hX3YJf+2QZe2RTMYVCNPCJDlVzVl1k
S86FU0JeJV/T/94gJkRgsxxfI62j9oR9//W7aOry9nvfveC8LDPg4OFD8gQQnQYj
RbOIVeZTXCUT5cjG3kZPksx0gkfY7ReUmDV0YEJXAlPrwkoaSzBj4Wb5zj6ksP59
GzL8PmR634KsQ7CVSfKDHIi8xfX1VIapu0h5O7n5wrYJQRnDKRT6EQW+0YXaJJnJ
IzGUjyxxH8/5cRtfyLp9wKTLQJvOmKohmYR94QtoB9esFNVaUoBoLtafI5LcNZe3
/x+QWDNlVJBoqbS+xZgFCUrwHu8kfvsCvGnVOU7vtFg4cbGEFH2Y8ZXyEsyj3nre
wwAD/w0E57aPfwNhLQbGlF5XZVsUmfVltTnfeEOAbJ8QNdQNJG6FZCZcAHYtdZbN
scUH7m3gcCjd56/jEPrBKmGi0TlpFFo0XqnWaqBxKHweJBxBqxl6PFZ9GSX7mWwO
yvZSOp1D+l8W38Z4nAPH34VX9dqIWNQ+uFEiVmat4y8tbVh2vWM5qn3Dv9eM1plP
AyS0a55e4Z5pf0SSaun7KlUKLBcqiSPDzbr+clGU0InoNk2QScq4D+C+s4IuaY8w
IjpT1dmAabPzPGFLKMALHCGr3nGU8lAkIB7e6WR+3PadAmCfaRduJ948whDusdNW
C6OqJnaWKzUpc7QNjB49ezsSUWSlwUkg05JX3I0rP3cH4dXEFuWGm+XaKu4gItxC
5KV/iOC3TfkeK3BJYtbYZNtL24vtPk/rN+8QRGivIFUpHyU/WcejdQ84JRq1IIog
I5Je8K1MU9Y+UXJ+z6OWGCD11hlxl0EcIXsV06wL66XoER2llcV7pPHrMPYBS6cK
BT/2wVr3nMcDiV+hqJ9IBQiBONKbJymhvc5GY4RoWBc47ptUcOEi0XQPf1ytJgL3
lhXD8oAcaBhvrIFvUOXvaPecixS0m8LgJrGWRIF3CXMiJH2hRN4OXDrpl+uOme2Y
WazUlnvxi8LTxMd91UisdXZ2J/2dlhPO7Mm5BZfD2FbTMy6c5qyFlmk3m6dwDEGm
M4W8hTO3kADE8moD+7BUNSML7Uv9iDe1MyZiSpz1Q318s0m7yl7UV/5ijOfUyd98
ukoIHLoATwEV7v1LcS7smW+APTj5Skd8ZOM4lKgychCyYxSMW4QJOqbw++8ClXxs
GpuTzhheeK+2yV0N0nBG4qN1IPjJEAQy6XDm5LaqtwgZvBdrP9r7/YtiJIz12qoR
2FCgX7y9H0dkF7QXZFKoXJZtb7NUtbQJzV5QFNVttsemmHVLGzxpX48qo8xrTIPJ
1tmvY1XJS2q3645eATMJMCoDanzikj8pmHOsHrMfSWN3gMubCly5scSmEGQF1m7B
EmYdMF7TiAUHqyOTp95mdaSoCGb55Z7xXKohe/T/BrsOMzT9qXC0aZGAfVE+La34
kymkIowgRJJKJgKn40BCezchqg9IGon3bBXkDLoWpfq6nPCsPb8ojPrOzjQJ75pb
Ho4IzKchbuO35fwYp6wfq7fr3pW49coZ/rYVA5M55R0wWGNqv4LDB8fwJ6UoVEzn
Pvww2/TNx7Jn0vvC6I2KpAw9HXb07UMzpL3IHsaIygE8HoxLeM5ye4qMetoi9Io/
5VgkPWeDVlogFxwjPnKwBm66x6O4+nK7KaSJW116kCV5TMdoCnm75j7XMuv6LJtu
VeEnM0HOA3mWNJo5R/RZOuwThBQcubkQYoy8PbDhiFW9u2G/YrcQGYc2US04/z2O
+fDKV+oayu+OQjV1UfoGmxoRJXqflpIePAjEyQw0KwcxpD4/NRyyS4cmYMQnu0oZ
sbIg5NQoR4PzOP909kngR2uYPEk+aDxDB8EXa2wYTmvufcRq2AcuWReC3DEdfPsp
gbfEvx04+pEVmrXUsm/CNnop7b2iw3wq7sA2zg830Q1FTEDBNwBDpfKvS2JrdO0V
gkHir2v+DUcE9KEaAiTUySgA6lzfKJ9eeEYobiUA1ajrXqJBpa0ZyAOLeEnhg0lb
xpbmn/bqZZDBKH93d25jAOTqgSYV0PdiLxDGfFVOx3vNQ2D46aYG27EoHg6Z++UW
/ab5usSPBWFkb/XUYWXD1Zq1VqtLJlKA6JFjn4y8atTgs5bx6bg1FAbi+IN1oWKe
+tzGRKxAqnnW+9RbNgY9wZlOy2LgJWSV1dRQcRXFv1DPjCArCmpgKC/Txd2gapDM
YyvqUoOe6xc/hKkVcEGYauY6AuVeOsVmvC1q2f1N0rfbf8iJg+r8kNh1Cc/Aj47A
C0BSba4Wb/331vfLJgbVTIeQDLumn+qcDzCpvwjJf9RnK3tN67HgTI225eXlViHd
YAhXUYoiigWztS74n+BeJFOANUlZHN0mxfa1RoVJB7fVNelA3GumfJhUAOa7BBKi
cIBLjJXv7C1LTwFFvf2+jBA/W1dDmcigvSJV5+eW4o/dFGPZb+9qKF7Nm1IHyAgq
hUhJ0jAdDZjTcNKvx0AxKWV/qPq8My37Xhci85C27YaQD69tvicIHBQ7D13LwTzx
h9oaxBW4vLcOKxVlsG8Nxw==
`pragma protect end_protected
