// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
siQeDDD2mbq6OWfIo6LjUzGVzlhbmogGf2tc3s1JPfYUAk2mVceAE84ng1B88swFTtNZMa6Ogl8n
jWkqryHKssVMfrckOiNsf6tQdKDGqTEMV9V5Fl3sjEy4ihugG7ecf9FGclx3JR3tfiFgXP50kLRi
IyNImNFsjWdLX/oFQ9mL0JNhaw58GfxLeSWDZrK8rt7LEDCWYPRwKhExaRrcPoPe1aWOayiqdcuf
HhJJp6+iyEyLI9TzGupT47Zm+GEXxlW/aIFylk9aUzrp1ZNjUYe667CTfilrAci4S2+Ndh6Mix4A
eh6m1DYgfvh2Jtnv0Rj+asvTjhYngVe46VNeUg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 37840)
d7+uX98a8Z8Uc52T7pRckasDjXpuxrSrjXZ5Ens1TrM7XpgDcenNMR/D744+1MrQUPsKiSIxawJ0
ciD4dYnoy2CwBfRgPulmKdELi9CWNVVGWayNC9pqF6d9X3aPeznmciDrw0CuceBJFXFM6WUW1yTZ
6X/hvtpvX+6k33TqbkLKWzfoCVzH2GH/Gig1wngy5OZLH7a9mNZ8u2lFBUllshntWMIrDV0CVGYK
twN1fszxDg0bGWmSWeCskIVUwCnT8mm6z2HwPMxcKPC+Cg84k2h1iv8KTEGSGbmXdOJqCzppOuiH
iat9+EilWvOGErc3RP2bPgcr5F3oN7FQGd+QKi2C4TPt9N56DP5oyMSNCZq4vG16DFoDmW3NQkke
0gxV9Rg3Hd0xNTVZCWaBCvniwRNNggjw0uuOjZJ+vvlzHwEMWshyER2RTMytqIyc302YkCEM7zNT
b4LqV03JJpSx6wEyaMnt6nk7N2URk0LAgP+tP1nqtDLq9YzrXE7im2eLEurqzs40NJh9qOjNJQ7J
aZQKD5pE3T7G74md8eJeNrZWIUGd/14rs92heYKpqPSljMFXNs/cbGLn9Oa5QvUnbnGsvGxWyRzs
e89JauAvIZQINglMtjwzfvo91n96koBYr6epp7T6SJnSrSJ72cYliSb0kRCDpheh23oYQwvMUzzU
V0bp5X9LLVZjtT9qPxk4zbe29HTWP5vktYktM8BljvnB8PorSRWwCoiTGyG45ajXDz4ZIGHAzszv
eITM/Xbv5LMNzknahOqGGV0z57giexgpWwgVZGLWtBH++ce808ZyzEuHhaUBHn6jXcdday2P2PkA
ksnQkEFtZRxqXf/Xzli5ENBhzIU1fC7FN/iksjp8nPX0R0brGL4xOTRDy+hp7dDKfk4Q4BBa72ig
S2cJVgtnRSugfBOZYNfdCHTH2t3TNM4GNUWtvtM735aVe8C3T7LMNO5m3t2pUKRorw6XWrmmN/xP
Ntbu9COJet01/vqTUkonSqtubg95O2dkZOXDFH5WiVb69cqJrRGrSy5o2ISkEyufNS10EytgPhOn
qUZbeK13vhlei9pvRtZlevf7kgjL7KKj4P4xcF29kGXvevwD03RhIG1XzW4GaSms0DNlV6GfoLei
mkCnSUfdaxolT3Z8B95pTV1Zd9BaiJNe8vtXE9sfsQF8BbTQzZScFb6KGqKd+xVui+hZrfZJTGTH
G+hjyzqdCKmzAyO8lFdfOoO4fBfOfz2LcwultieALmd0VTW/9GsKzw8fIYv5HLHh9JmZpdadRBtt
ARz9FqP+MF1pHzEXJ5I8bWe55x8VDEjTHIFUtXBb9BSWfm284UcGotbmhXtj2Q5Ne2XnnuMDnZpn
1rN20nQJCQIwgH1PZib2CvC0cWXodzjZYahP1Bo+rdO2fTHE00FsEr7vSMSHiasylonMlRyMkZlA
Ahntn0CAZW9Kk3xm91yqbKG9DPh6DodHMazRqVAu0O7orLSiRjPerMj8dYGXzW3ZdciogwkegUUt
E0YLRL3bvp93Rr10GgjVQ/0FEmci9cGSazaVBKIU+ilYlXnTTUQghM26l8qkXeH67xBvl0lWN6Mk
PrpS4sp6Y1ywJmQGdjDQghNnuWHTSm6jkoimwQoKqLcEmfiSkiZQfRlz6xIdhQP6aQXpV70jnd/9
Uqkcnw5uL1rLz6WeGiXsqDYBHA6+v/a/m780jViYKu4vKZ9xTwg4Lrm0s28gmgLzoBC1OQZ1GmAX
z3U+JQPoxiX+YEpLPA5ezbVPjXfUyLlfq5hzEahflOarbh1Bqg74RGUER30Ej2o3E+ubJ5BgU9LP
KeHgrNeeZo/uBL7YorVancAAd/ayFp/t8GNeKSMyG1YEdgMg5YN1xCh42mmameCReRFqobZCL5HJ
E1B5RrjB9EHPlVqWQfi+/4oyvl/sbaewQFKc9VBLDu9C5dkYoSVLUjLklMd6s1u6nph5fRzSPfCM
RRHCBOCaiKJtK+4CSKtv+mqIDygw5I5mGzEcfnw2EkeyucRg/So8+E7fIm1dRzbsc56xbsnEBYz/
zG9weFkQgJjTWtqGzjRUKdWp7zFyx3MHMErfFkfI6J3THTyY20Pa43n7aEL6TsdVA9liZsh58kcB
omrgZVJEKq1a5Ie9hj+yPmO+X3DU8gC/JiAm77z4NaK6pgf7F7HVJg4XYkOV4cb75WPG5kPRYDK2
wWPo49jVqWdCxWYtvBdHcy4AhXlThEW4yUFMirl9iykqRWRSh1oj3nTuExOYc25j/iAcigQq5huV
DPR/xNGSwCPMhkATnafhT3RE0p8dWweFqsmO8QP22HXZlNqaRlH6ho4AqCTiQzcoLtSijvH5U2T3
B8RrtvzJPXxoLYDFlI8st603lQQdzi+gEDr2xaCiARDcNmgfWj9H2BIGEDaItFsmy9SBLubtawOp
lUrplw1zN4CmCYo/X74dtSWezMW/oyfvld4nFS++RQ7zK/MqB1g21ugcoAPWX5G1u8jKMFQxiCHb
wa+eNEZCGXq77oaMIBV2PR0Iwcio6m9c4ictZcV4jFDNtI6ykbIvJq2MmBjVcPR6HAzZ/XRLq3li
Nuzh0DIfcMipv95lX/3RC9y6cIY2jB4Q465jxPu6eeuLTHucqYYdzcGFGbwEmmrXpCP1vis5fqSI
IITcSVcLUFtjUxfdodUf/KfrQ0gx6E7mAnZ1JiNr9gQhUF5Ngj1lqfRNlJpxHYfQOUPTYSMVjOnV
JpFYf5YMQjZpR+exrS3Z2udoSyKi/Z2VSyst1gqOY/URdJcYpUoma7jfuOR0V79nOgQ/NKY7WBiJ
ecHWNW2IwsucXFkE4bYqjtwpPWYW3OI7x5rNafs7GEFeZNFygfRiUitIWgpdrLnnlTwTnTCvNdBv
81/lyv8Pi3lF00+Ns25u9FQGP2SVhICsxxfmDGlko7Y4QLXADSMc7zSCThKnEaBFtwh71pIMRDwl
mVH5irdxw7AT6t8Z4WKa/7WHAxjaQSK+6t28Y+bLHavV8Qw+tKU7ACFXbvtyZwBqqP4vSxwB65j5
z6C7hoPMWev032v7eRDH6Fp7Fp3hox95SOyLbCR8TVwco0a1hcqW0xQ+r5uhFwbt3Knez+xBmvPp
Zpt3XGqRsQ1uz9Cj08eUF0rH25k11KeBGXsXmYfd8b8BVtB6MVPOuVmMjfFV7RzeeL804/9fgHdS
8VjYhQsSYX5U0pfWeFSQPfapvB3poyJDLPQMtUUspdVHbVtVymo/oVSvmmKOH1hX2ko+wY08oyFo
afsrVLP6//L8KYdIKcdPCc9Nq71h9UgZ38tzDivNFKMFFI9sfzdc1t1ZhKsY79gVXs4oFvDEW1q6
Zby7+zEkYZHDmYerAX93C1lEBN3r6k8axRICHSOMfAdXPmkYnPSs3qHbKl0fa0MY4532ZPkQO4tb
rOIJ/0eIR3JLVYDjJOa2p3/CzJIBIy2ktx6nZrwBLTJl32u12kGVwjCABq+xGWC/AOj9vY5Ga2S6
UkdDeIVkfiw+sx+AdyHyYAKIgzXMfboOAX683lcDZ8eHhVVnAHk4ap80St90aac+hhBYEFODiRU1
R020v81nN4qlLKCcIFZf34CD0NlkHYolY9OShVtP7m+0po71VaUFGVDmCMgnLENz4IKV9RFWyM3M
ZoE7tGJtp74BxY+pX2fCRnlqHTMKadvtRkaMtR9STTQlKU1OATAHFNpq8vAh6RxvTFSchprT2wu4
V4Xfk7pc1sT51nqqTBnTiz1W7LN01HlekfkCaNNJamdN5Hmxpyxw/UVYcxHZlSpSoISE2hki7knG
nx6MOfUW0jizSQSVEnuU60NqUHfIfeCONpueZ0oEQ6rT7s/7wYAiXLdFOe+q/GUFNmtRd5fRsmEa
hH99W0xnO3TSIf6EIBxm7TbUCJGN8rvd0C0ZwuP2JaXR+x6uyLGYCPer5Te2LXNMJpITj5CNG5HZ
4/BDbl6lWARbwRLgGeffvrTrb/2kzurEM90lDXhFgqQm0af6gTonafn+sL5ju4o5csJoZ9ZROof7
a7v1Kw0kDOQoM1hcU8C1Fp0kEbLrWtNbRVCs+zQfotI7imaI06CovGVZ5GUcu62dyQj/tlqUzHMA
MrQgDLHGCnJKAUBlV8MHodGTHocaqtkrikkgXqhGvlMi+c2yJrxyf9uLzHH1rPA1mO26PeyZSJlj
MQAN5z2u1A2OXGlH7J35C6I1oOzFkbICLkcn8uG4Dt5/W41SEibP50hfT0D9//+OZb32kSESg2Am
pwQC9tqZAksTSgsZ1Y8vzYWLK7HjnxB5ODflsryCGfGJZhQbCP43Hftiz0iLPjtWCSZEIplrf+w/
UZISQBLvsAkvjoDVerT6m4uCancpIC5GO+VmCNlpvjuEzXOzJ0U+Z/gFSMl7FUcCzNfOBkp0AKNQ
Fe8emxZydjI5ysWVJHQpmrfqfYU5CXoAde8W2mDBbM8bexB19UVJYjpZzqOaGI3OPq/kYdGPCn2a
DHJNQdkIhOUvPEG8FFaoh9M+88OIvZr8+tEcwzFjFwbqt8YG5q7nUgPiI8VZUUZGenruo5AbQrBO
lMiK0iJ1ZYhEfjtn8yTwYjhJK05RxE/fydovtMeDHErm5kKl3aqUKbA03WoNzMjoRmQghvChu/lq
pfa2VA0HQXs3RO2j6Vl48m0PD2zDMy+/0uuJBSs85jQlrMxFW6xgTLtgvbSGVT2QU2fPmyLUmmVq
W7dwdLt/AmrLcTpkFJipaNXrSf3uOHzcBFkV4ga0pHXDdAk6WKjXVyWy5nLjuAzkT/pGwJCfmPWX
XC7C8pMttyoP2jfiKGVTvz+2H4hBKWisrGkZq2bfieGzLpRf1GfWC5NljE/mpfgXRF3X9i3MCAsG
oodpgXX3LwSQsmMsQf5/WVIs+VcldUvjNN6j4txCnOLehkt9bGF7xc32QbJ9MAZod1Fk0FFMRMMC
z8MNMjPSebBA3B0BKO4aMLeNCcuE77JdQfPAlgDLQgG3YR94lQjPmq5+DRnf19zESH4tFOlmBC7Z
kO3/BM1a37iGuKkTU14C6MfomU4gzkVdW+YlI4e6UeidZgVKVwxc+pnepYkVN9roB5ICuEKYWa+2
ox83WJgVe6Qbio9cMnzP2nDg77s4e4UyqaY8kZvVXnYntbN8oVc02sjBY7i30fgsRuKsYtKXkcFp
uZLc+Ksm42Eb5VzUsypBQrqMrTPzj6DHJwjqcZH8HeYHzgpjRo8ZL8ZYKjLn2hZoTuhHxCq4Rv1x
r04HdzZLzFJrXgUirlz2DgpBtEWCQrPaPNcVBPPKP2m6nU1xmuDIjZMdgr4nKTpuviiOkUGg1rGL
R0CSlHsJ6DfUUtSpFe9284nuTWARSrtShn2DNGcM2nXElyHjPUmMql9s2zBum3W/oJ6s1TdqnoZ6
t41eZ7WfnVUkJieRmNVBT3Mj1RW10TQX6MeB91u4as3T7WAyum1HBEVkvw+qnKVq4mwtBhgksI5W
UqjwPhPFUvYUaHEEtuN6B7MgCt7WH8FcvV0vnwB/vsziJEgd9iihvbal7AufswSDwLgXQCFUChM6
kEU6lT+p0yR5PpKLrB9LyY5+cyKhXwelUaY94rWtAp2DYx/qlHSGqVyDbQBz2xFGFvA4jNbEPolL
rmBve/rMhGH4VgSfuKG7WZWd+qB3kMNePUkguoLqdGOm+Ywl6clYD7tEup8DuoPPWXup3lRVUTPj
qnZnmzbNKY9g+mXiweMrz0spz680Ein7CnzBx9eqKDKcf5MnOtgYu23lGDCDKEFy4U1yOTeQbC4T
U61qAxH2Fn3W1SBfZSNk3mAhSEund1nr6nm5Tz4TRqIPnKwQnSBpvifRBnqX36gEMP/q4bxqdINp
hI1B9cIWWqaY+Ezy4WNkNy8E6lEi2m3fJlGbxy/musZR1HQBa42n2kR23Yg6/8YL7kbxQxJxXOgs
b/z6/+DhkrMAZZ2f0DiTxE/VXddBqtuPyZLK/rcK+QrD14/3R8BPkIY7hIEIPC/DtaGty1KhfMi4
bsygyvWnVIl6MBP0FGDqtNAen5Uujz2h1Hnbe0k7hc2Jh45bztmg24YJ9tg8JoGf7bOuqEo97Qy/
4m+Fr7GcJJSaWTxF6BWHGspz6bYLRmGRjExz09e+SuoP3j6Ns7xbSIqa/BiusDQXGlu7Dod7/KbM
LMUpcfjHmn8T+L2lN9Q/t6FA+EZx5un96QrTNug1zP9yOScIZvjCaXH5Q3r96eUvhBCZHPvG8MOr
6Ge8rPGsGKCjAD8J9q4HiKx7nj3ccUyUhPzjnlLRUmF2XEbxtdaFr6MLqpJSxs40Lny0HwwQHpIT
24qO7CRvK001yAhSXetizUXH4v8as32YC93rZw/oZTE+fl/YY/z8BZcB6OcH5l0D3Zt4DXrDPrOy
rLcYyZ9ASGVgKcZaGWndFffAz0ovkyht3Yx9WzvqPxp09xwekgEKbS8qurbwMic+QBf902yw9N57
F1rVcZ+sFvwI3XYfS1ZVSjjsGrIErhHvoISV0lgA0W87h9CHOeA3e+4s0BX/Jxt1EPFozTZJSLZ1
xFiq53lRDPiBTCdwJJglZYgIZoDrZd79DFDsLD45FJunwjMRfmEHCkusb0Qn/wCLnNw6p+YHAdIC
2hLOubzfd8lxhdPbJX/Kub+oroUXCaBcCIEQTB6egrWz0KctdrXFO0a6znyE2G0N57FF3u89VmKK
nUnuZxPyky9KuaIplMXwhAbHMP92B2KmOo7aodZ+UVhLeVWa8cBrB6/3n546YWEcK5BVH7U8q0Kw
cjAqWwnZK/B5NlkJKriVjSX/SlP/3quicw5vQYAqszgCpTN/Re7zEfbybpmmIU5s/2m/zsAtAZw5
JcITXpHCeIFfSnUR3hjlKD0WM3xoFnOASf6/XGKPmKv2Ds4RISp1WTH5FVG3NN+JoGJrQhZlJtsT
he8nScKFzZuDklE1NcUiu+1RH1NBltIspl1tmr3t4jYZvkZ2+kOu7uD9/GHdQ0zi9SxVrmggFffz
IsfjHqkjZ+K8I7Coj/WcJ6VDEmOxhQFU9Etr4VuBlMSfyWdWyIfu0wbtCorAtowEvk7S5fmjuGm0
Y+DqLXPSMgcZuljKl6Z/OyMVgKXFf1fnFAeDxL0OxJq3hdSExPkj7dpgwQHdXzKIthjc5hAPj5jq
cCqU7JoOn+dnirqRgyjEK+MlB3l/s+8VO285K4u+5nb6sDxptzxkvygu6v5wfzxCaURC2U7wfcjI
v2lv2PHUxGaIht3/5NsPpss4Su03IP0GwMJaTVT5hUzC7YsTQfFruSOCmdYs1NNZjpEP1zX7zz56
kg2YpGHyTESw0M8rgWIOlZC6z4YCjq78ZGjaKDhV216qWo8ywuPiH2jOs7wSPakX8P50QAA4LXkv
BySRIuOCjZ40MEMjJ4USXk/11jE6vcu7FdcxAuwVdUWd06wbeMCeKWynnIUJgaqFUY0Ri8wjbjEs
bd4YSc9kYYhqfBi+7py18DfC/85M4wkO+sKrWSn0K4S6Ofzob6f/POvFT341JQEwhZtPi6MIVYmt
/5osdHfZrJNZ5L/A/WTfXXCoEaSQB34EnadwMDGbYrvCZ15YdvW4KuAYH8kqfHq+Y23Wl1YZ0suO
jxwlmPpbrGbdlcH0MiE/JcPGA+BsARkO2TY+4b8mWrbrMKb0qLEkHPjtsFcMfirD0IRDrZFAdgcL
RTpm3lL5QraHLnNStVWJry/63o5txciGEID8jmuwhTYPbx0fiucOAcHfr/j3wTmOnCbDJZxtRq5w
VMWnBmT/KGiQXLxMH3+C90zllS/s3rM0MAc3PsmCE4dWm0MRnPo1nZCwk3EzrOkao/lvAHmBGl6p
KKqUhN1iL5v2JCMUfJzQFIaGYsaf68vqpLQ49wDI9nz4F6ZCX+gWv9Bw1MvOY/w+hx/JaTfREM7v
2eJ7TJMWEgFzsUkdCRSxcEmGvVWtHGB+54WAsEaJQVOvzhLJD1ddjFqag68pyeH8rPbKBD5ky/wl
gZX7Lt9AVrY88NWJoswEpSgz/dDmdiexoZpgeYB+1T04Mde2mVCoTcEXJo1/rx5XDGF3JlJBWXTD
KUG5yTubEvCRyXHBZmxKLCtG5iZBkGIpVW4oF8GkXtErm8GuxpqR1jjNJeeHNH9+zTTuHpnDVrQ9
2ZBk74i+TNowK4Ntx0jufznKEfdRPL+qYJMLm4d2OF2RXXzfQWa6TyDQrR1x8m5U/4bpqF4fXOq9
s2pKMeMds7KWcMERx/mejlZvsR80V6OAC+CYM8BzZy6tHvhDwOI9vrtslCFojjkB6NyzNo5Kp4Gi
CbrrqqqmwCMhH+1WFiEesf+t80Ko+KpH+tz5mY/KOT/OV+/tfAT2eQJxVVa6MiLzfx+nPj9FV+3l
WjGsaEplACnJUlcDCTZVlx3IbOvPOZlAqB6HMayeqZzKHK4VpxlC5IleK2AOIaQslYHagrhefqd1
sRwDzslbI2HccjPl0Buf8qFsVn/WzJKSs0/iwgDHYvW7bvfG04SG0tXGBwSmxMCFHeZQO/+Rrw10
nxBu0aUd2ALdsueDT1iW9lwOTJALQqXN6zURSegMXq+/vZId6oTEAz3LS72omNP5fdelpHTv9ve3
Jhar5m+i6S1qL0BbEPu2s/1wa5ENCNBoY317dbLZfZOYHQMa9oP6IPM5Ce6pnLs8zeCiBSe9Iw+m
7miWs8cYXcuHuV9701kWtDE7Ef/yuYOt6WHQ/J1sSPdBhKOPWaNTRgPVDYKnsykLkyrNzlIJojCT
2273R+juowzW2rgJXmNETXBKhHcanS/8taDYskuiQJsG3QtHUFCKBVWkFrZJI4ZzoNxbrQhEuJNJ
3Dzr0SO4/GI9jdnFpjuV9sCv4lcEz/1zNJzzca7nwaeIZEh4+ZtnJnYAZZ3tqRfZ1kiujRM9d4T2
FdNP/PEK/8aiUPhla715THNg0GkUlppss7ToxepvIR5VkWf36QWQlSshj7uwi+tbEEEy4AwmJf4+
3QVqRZRpPKoM18MBhH10My9geIhyuhEYikQ2WP3w7AzuOlNbE1GDLHZ+wPogMDUx2e9NdvaqYW8x
eG/SEv0JkU+PCm+CW4oK2MHLkoA9qAWaIO4YeqtuVasyQY/jX54HXHQ1HXEet/eQwkW0sopDIyyy
VxzU8r9f/3ptdxyGApNQbthiF0dH1aJOigtDlg+f3+TGEq6fgKU/q9DVrG3VKxhxG/dUp8bFmcnF
2eQNHSvhKSwY9sWvMGxEYhGoRnK5vjmNp9v+dIjHPg/6vvhRFhTZFQWedN/GfRa2AK8k6EhZiQKM
dsbmppFYda8IUCq3l7hCZJFD9C/ctG19tGh+1tVvkuQg1czy3cZ1BPgjNGzZ5fbKosNJol3W8r3J
kXSNQnrlv8kHH4K+rSQI8nbYIgFG7NBWqJyUU7vTFhec0tINMgLnLe37DbPA44FsxxIUI2sl/hUF
Aj3g3tFKyLXOCsTgDjVMTVjXmgFUQVUUuGUJdOQDBWglju8jVLGRhMyBbC1ylZ7Ik0ZdbBd3OcsC
Ua3DBZtCO5qsIEBNtJj2dPUSJBB1Oy5/5A1mOhwsXaVWL1AE153WEFg2e/8CPHA+B18cL5uqLFIQ
/S/N/SiwKvNA1FGOAPxD8Bnzm8EvQKUNpEffIovDVTlIoW3LlVMOWjegWPmf1DIr/N/DlYXh59b6
lcK0PT9nCEYsx0UyllF+XnUIwkpIcdpY/DcfLtdIAu8fZFRtCLDXPaDdxDuUJf2tbxw1iwkTLcwL
vKzs8BDFkcY91MncCdoev8QUDrx/cHPaonUr/ZhS4tltEHgFOcrsCRaw2U6kRyDZYVooY6p5u/mB
5thu+5U8d4HJOhSp/fdmw0tJx3hDmFurR8Xm4aDsXKCfONu2oqNbsvhQtbmkU/trpVQ86Yg0HJ8U
uC+9zB8bAC/pnudVsYu7kFFhwT8AMZIqb4uUwAUyFlvMIPQKOwU5g2Ooz5FvkB4tEzaN2wiiaWcY
xNgGpJRieCldLlfUjMsKM4aBtgCiolEbswjg2CyxVkXWGA/CeUszqp7zfIIa0zveL8D8COj2emmj
opFzPfq/EmRiXar+/RkLomLyYW9sTA/hZds6M5kaYLMQ1U8blgxZObooWlXzym5kcgEvDwzqR5rv
qFhDdevPCPIrpqhtkgVzVeiqIS9BNs8t5OQDJzecGx+OMWs53uso8xUorWGrDor/1ruwycGj5nLp
ZZctC2YZEkpIaSZSM02enIpPMacARrIDhN7R+GuYmp+9QJkqw1lo1G/KFRBg9q/uqCBr4VkmGHwz
CtpK+/XcuSg4UOHISs9fk9z9J9Kq1ZVK5bMHJP2ojEmFDSVtMPYR4WFveiPAAPCVTTgxYUXpaQxv
oazV3j0/Q/vPPIqtEReCV5jJ6B/6pkcQzh+d2fiSQsOMwltsOYP6XAEuttsGlznQCo34aBiQZ7v9
CPLQ1K1oF6eS0z9Pwn7IDNvXtUWkItzyn4AcQmGBVxuIQL6mKBUpNPxzYREJ09DHcYHS8iAF1fQl
Z3Vh61JllPxUyASDZMMI6abs4IbPudiVs3Ec52oLjIVsM9AZDcaa+eODEQjYWux1tBOoswPYEFNp
2qsqwziHMpZ/gAYceLQ+FsXjQAscAwyrO5S76cKCmEUUnltgyoO0hmKUaupwwxgq7TjNDos7qISA
/69MRbXT32GF54RvbHfAvCWyxkCXpSYST+HiyrgGacbQNncdG1t2d8AZI5mCqe8JgsuLHXDVJF2j
g1kYjf7IimBbf6sujBPLj3cYQluGhwgu0sJZt0kpim1rIQqZB/p8UEZVfeta/fPALpUScT6XQlL7
WZ+p5wrjPkDSSUwaDaQRZ99TvZKbmIb4YBVWzVZhcUTlO0nLyNOHto31G8Z6gjmK0+FP5cNMMgaN
5wANB7DQTWKTsFJQTMxYU4FAV/aYGU3IlPuBMFb0IFjok/Pk8AnlIT+TngJWiIU+Es83BFF6W6OJ
luh6HXpOMNaXk4QiY6682RONGaAA9qdhgCSORjd8QiPwv1wJ3g+dyt4SLpkc6yBg7qd6IfkMQkj2
Lhr8XwY7FZ/P7NIB64tsr8vqk+6TPBBQGOqKpFNfxNI1uQV/L1F7p+4X11cdWNW4QdTKv1CpS8zG
1PrwKEFyWpODuDzLmARK2/Ptl5ZzvYgugeRdm5wD1kISWJuiYhjNPhrPwo+1XUqeeJNFshhSrAvD
n0GlFyZESWngE0as/1L0nZZ7fnq9dtLNMfirCB44lOXYhyBPQ0cbwiHA0QajltmHSuBC4HPV+T9C
JNcbFADCXbVePPUMyCv8seD6AX76McZXdFtIwK9HdjqFzhcRl5nuw04CzGgJuoiGfbHTSMoOhBn5
hpj42/dJAeEiY2uKf9MNFGZS7qfCWYkaxHZ8s39iPuKR1Rf8M27UlbJfN8F5OjPAx28c3YJZXIAs
YpdO/PLGq7tVwxcq1vJNF2eKbwvUb3hTuS0H5PH9l+F5bnWj9mPX32j4CnPh6Fd3DLNDyRKNhSZP
98VMD0v2gGkUBeGIEtnTsnAEbE57RFep3wNTQt8GwAj1o/UtpQdhOQUh/EtaLEGg8YCNG3RrYbl1
gERtXfzcWhfDKHeFiHcHq9eSAIOhALCaROCPLFcAKVbzLkXC5OQQK0/PBwDdDt3sy7r6uI405QB4
fvSLjDKBYFwv4yWw6DwQrecS4No2bk4O5bxplWY6XdeP8SrRjDYQlCPpq+QFkHP6mMdPTqfn1UJ1
jw9xLxnsRFZxg5ehXqDhtz00pJZvfAzjSSiBPXbB8RrmnoW177Jak3N8A6lXUTK5i5YcYNW0gecY
CqZ+gQw/veiFVRvEpbkaliOLxCexm7xtHA9kxynSGN03hTvSqMsrL7HydR/GeIHq2rlzVphpp+Zb
ITBUSyKdgsxS8e5qel6PqqwtIhnpGa7mcp0b+/FyWGZRgsbaiSvj54yzj2MEsQI5ibXbW+TtYS3J
5ZeeTRcZZDCv7TGnc7tGLfp5PLbDMxIN9ELiycAarwFKn7WXIq+aHdgTwT7E7wQfo1qBxcPruOKe
WqfS4D8Eq1zx4PdqaTfh/tnR3Q/xeQ43eDPOZkJ0DOvZYoFm7g9BJKE97laQ6EaddkO2IgQH98S6
0FBGfpdNVD60oLAdaJJh6WREFg90YJ8d4EcjIEZ4et1ehYWCaUVV7qDWclXqaTvvBt0DpiAzjwY9
b/NKDGk29lu7I1/wkfITsjP6OB5j5BzMoqpwgbyFBLEM+37hLWS04TePlY8ZAOXeuN3zMRXpTlBc
Y2iTdrutiHOJmZs/4P+7u2oxYMpVAucrg5jPhWPWmCac8IAtf9trO2bi5d9sJwAOzQl+PFvtmY4T
AGOWWqwA/AlbP6c+rcwF8lKUXAm/Po/tsCQ1kmnSg5YaUHGofBN3gaqSr7Ebo5upIVY0CcxZJBRt
lVfbs8JY19stVhss3UHQ2XNN6b50HYvHjx9jAgXDYCmg79XsVDasYcCRvHYMp/bx2mWl20sRad/A
6Wqe8OnMm6u08xX2EB4Ar6x/JTeiZmuPORZ1FQ73D3gRPIOf5MUSoWMFhwpiMriSNlwyPq1Nn1Bd
8m6wbjdiLXK6JfOaeexB6K/QEmLovpZw8Xr+vhj/1AXo0GMCnBVo7Bk9vvEqF+J8yXkIjYGQgZr8
zDNtEVML4YnfcA3piS1nXdXyGb3fXiZs83R1W10iuFeeHakHtzkzbQA/A/Lf46TeY/JqPyzNmEj9
lKczDBaS9qnRI2Tc9kbbVSNThqbCxrwjtzTNpRr/NzPrqP0C2h+UIya2SXNbAXwsLB9+FSztt/mT
n6MtsBzEj52GAlTfYtgGarUSX/s8ED4X1ellWq/0CGQUL6AGjknwqbqG3jvOSuoUj0amRPxo8d5u
QzYupXqQOHS9mPXSX/gDVPkaNJjLHqiOt7PDTX+1eYFYRHXP5BxsLstf2FQObE8mGcaCqmPBBrzm
h86mPk10NYxQJ9XookOJD4ejnded+hRk2TS6R1+A9kNe6kB5003/SYRAYl/CmkbVKcPI0uJKLUjV
iRgmHt4i4YYlqL8g+xH+doRdhNxHXl0z0F26mVASSyyEG3NboQLwHBfEUyw8mXNyvgVSgSCBCjBO
iVf/VfR/BdJVdg+DS+7t2L7jCTSCoptgvSnIb0u9B2+Hmi3KPUYZ2uvO4s5bHIAWBFIpTpWAzxuB
FZhf5P+HMIRiUSE79NZBZjdAin4BbzBJ+IDgvvjJp/fBrDFQczPmi4OoqTXWxDBVGAmle9yg4Kl3
3Ut9KzefvzMWADO3mjjfK52jmx/kNiuai6NfSUiYZoTT0Nkr6QzXVYTVxglzW80uyJdP9Ic2jEo6
k4AlB52Tt/kVqvxf5TnOkwQI4m0e6uRgKb917vD+bRUpE2Ycfz1i9t18s+jpM79uBlQbbc4Ay4TN
iVtkVvit8jYKJUFKFF68/PZ0dpS0StzCwkAs8z1iweIACflSqx4rUSMWi7rTdQ2b6Ae/WgNsCVsk
y/DGvCIzxLwbWKVP/qmBVa3WE3DnpRpsVxAv80+hZYXa+cWk7gapejW2iUcCKg6Ue4xuv1EJGU4V
ZSes7kyKhF+DtGQNBJeB1UyVdknnVeHcKDOVUAOnVVqnnD97EgJ6SzRmICh4YvHS3Ybhk6dx1md2
ztOr9A2G087BVgHpH10dz7aOo7pNtK1ET/L5WEhnta+Pknk2ZTG0CzKtuYgYzU7Zk+r5w8GFPR4X
pVrm6shxYtrhQWio0udAlEFRytm/cLnEL6vGKmPDZ8OxL8spVU3d7ty943d6xHFbAEa7RNW89ztC
bQxlK2c+sCIpBnq+R1dJI9gToQDMX3Gv6SqjjZnah0xiIq7oPw5pwP4K9iVN4+YU2tqwx++NzREj
Ke/3nDq/2Yj7GqJpsZyPoyZpw4GKBDiw7ExieWnr143ZtmsrJ58frIRgVa+vvAZT7yZ1KTMsdhaj
7rZznAu0Qk+Di4u/5HtSlMMEueVZjvoRXZCHJtIb5FJ3CyUUR44ExweEc5DcDHVWRUAA5rFCTwHl
aiI7OVwpG45OgFvKCkTTZUmtyLoNXziwzVXQ9+mNBjWfe2/z0LJvqppitPxgqlfexkXi0n6GF37y
fg6zpQqwfgMoiBxZoKiOPVLjzMihco2oMERjldbs6XFgThakJRbShnv3fteEHhgez2UjWW2DMUWY
i4yGSg8ahbde65LJtP6brfb58L+DlKSh4RhS//RGAvmwFEqCw9AMjkjKjZoFNyM+pjDVbYPC3LuA
RZpn24yXQ1aVDleI/bzpUM/y9G29DwoBIAPIi+W2Yi+NM6nJGfeKyYWpixHXSQga0Q/4BlL6PUpb
7uQV53zGdLvXAJz+FuV2uMySNxlikdCbbZWOYoSLHb/nBOnrfZ4LxW5ECGGeV+psmcw8+MDcdUhi
/bBB2RjnEduc+lw1CMMfcPBlCwerlLuBd8uJZ8LBNfNsfcOo3uo5dzk2RcEP/dFCe6xScAisKzSx
9Cf1yoNrmDql/yolbKwDNcDm0PnX7NBJ1mS0yRppGATXtLxrM5AbZmqMtnjjoiEWuKWZ07pNtyKw
/MxheXI5VpSXEr1Dvr/HkHoCBm+N+WNn+3NPzgVRqIu8sNlO8dStw2/8TqzF+lckLNKx8G7YYt8Z
tAbbiZphHAU0yZopVoLD50WXdlamYKCavv04CuaSMDvqVqErI0Qs4SpiQElTjnPV4dvofvwwoIW3
5NNOK4LTfd/RZVKxtvbXXqzOA5NVJavd8VG5y/tuMXCPTBQ2iOCY635VGr26O3afnXuJ/vH47MbQ
FVkzS/4WCzo10TqSWDDdWW4pm2FV+/T9k2ptAGmPDpO+83w4sP+gTsLj6a9WVjMN4vIHTFWQZzs+
MVnwWYcc2x+uLmcQXPEoXmssXuhxcpYiL80cJc+oeHJjhYWKXv38Ld9Dw5A8V7N/5vxGqn9jm2Yl
a345nY4K/8QweKYvbmhBuuUbj9R7mZWg6z9o29LCEPlQD1bb4WpH0w9Dw+8Q1ZTbQvOQugb/o3Wx
9mZEjxDj2LSr3DyliqizqqeHBn4QdNH8gr0DCzkQ6RwmecN7Y0/zDJYzBB2lnfgSc0xgEdB9wr+n
O4btIjWDlw8FcKWmn4hfXe2rRUD6oaKlunvkz7AyOHY6zdTDeh99qtJjcGdxnsuOxOVbJ4fH5Bp2
Yb0Wam3yrhSW0LbMi3QVDX3dRco8hDfg5RTjqMctSobw5I5TSmBxesTA/bObnrfpauWxuHKbvuaG
kfinh/CIlSeRdA8C3NpDJP2JobdSxqj2n2KQAiwCYVcjAB3DY2EHfrJ0P1xycvnkPzFRtVpDwUlV
pWL04pbNwLxuBCIhrgvJdjCBETEpfhUD7+S2DRGh0PJYsqNRvqb40PX453S7gw2nrXj5cZiiK2lH
+AveTewM5i6COsmN+3Gl9qGsjjAWqpwylLM39zsVhORhflf4SK1AkALBT+jDSZSnmALLeYOzguLP
qJGjtLlGYnFvlmRGMUoj5IuZ9NdP0UquPv7bhXEbCIBrnKId+gatmfvvVXLfMWdiL6y6DvDKFlhm
SQ4Ekwz5he/8/7lMosWxN1aaZydki3/d2paMPb2LOAUzgaUc7dGdhyMB0b3+uJFwt7icikFKfd2a
XDwx5lcQYK+NxtVZsYAkgBd1Dv/2lyHSEirbgh2dsS6FcTMnepFOzC85gINFoXDPvdCK/XEH5sFu
TiorDggXJVvduW8DOTv0adOr0fsE+FfrSaUjnGDU2XmKu4B0qkghOAvE+uBCaHji6E/5wec3lPa5
cyogokRxARxVyOn6T40oliQoU96QnNbnNN7c4zlLekUfqJVHV2MA+HUZPuOJSELUBLhFXmEW+dh8
hFZbUZndCkvpeUoIVaN1yBVtk5xB5nfv6JFLU/Zn57Slhu7UQPQ5gOGIABkjta/EOvuV6VHoFNmd
8E8aTBNPSvj82oJOGP2CQgN8eG0DXmp0XtXQ0tkvLdd+6helEUOiukVjR/2nFM8/xT7WAx25cD7m
PEh4jzjztbLbMNEGSY4Y2YPHNeMf19IYdGT1NHC8FV3qnJRwvS+p2lJ9IDqt8X/uxTwABMPk1rWi
nfRD2fgmoizf/EOKtA+hprxlSr8mM9h383DLjylO1t7tHoCMO0v0Jhq0gYorxUhL5UBC15yJP/8S
0Xa0GNFru2UH6UN00e8zXPYmHImBqnfq0l9bBzOB8WPe4fQwjOJuEC7+x+E+7+TsFv8S6q46oDI7
InmledVIl7ibOEp0i0znlBaJ2eIMuib9NhcVtOzTQBFAupYu7kEhRs8fzAOe75LhK7Salu0zlnTm
SdG92pNfgXartZNhKGC5jT+1aMsocnetGX/43RFhjF475IRUwrC3bxhpiK0rLwkKskuxJg+ROVsr
m+95S2cwBf/0vSrj93NMoiCQGpB2mS5fYiQZDSkXKQ4ESQ1nZ0lA6Gq5C+RZuL7isZzyYSJSm6j+
WUgavF4YY31pZXDqELmJGaLytENPIV+7qaEGiQuFCQhnfrdQo+eoMSZnYomM+eqPmf4Z0AhZ6I/B
ITzORLr9foA1ZoMMG7kPPuZo6xP0hWuJeF5qyh4/4K6qZoyhVHY3Vmn5D1uK8kpqpC2IZEJ80wYk
3NlSaIlp9I+3llbMtA9B2oT4f4hXOYHz5R8+Osxz5EaenJx6Ddw5wRjXWCBdcEyUlqZNtMgosg5w
fxPS1sMwlk3+BDRlcg/KZukcXjd6iifMooHico/HezHgVTY4rXFor9G1mk0r91N4wD1qYDU+2Uvn
MWSJr3tGW1ydd0ULax7g5RX6iPrTkysT4E9nTIyfKPHFOeLYAkERB7mih0KHwJjaYDvFyxRL4Gj2
ZjLIo/VAA/5ch+PfSQpga5VyU+oZYuUQD179SuUHv0hMO2Jwc9fioGME87LFYTXfvCTF+gTuqw/d
SPls9IJePOpMHmGYrKNNhrwktv3fHxcJHROCm4pHSnMvbjnvvLuAo4iMFdfkZAAlzUb6nA599o6c
FtckeM1qAVVbSj8339gD/IuFbvH4UTD8TCj8fvCjCm75bUo96wXs2jZixiW9dGyeRkdRON4CFjIT
/0Sfa5ru9bE2TgTIzf5sf6bx7Nvl8qdR1LAy8Ur3XK8963uqU9yystKgnx9fvVWo5ZeBuXN5beMv
AlbT1OQX9WSPoma11WKrrJQEP2BtZvsWIK/4Yv97tD+kshl50lMb0Hxie53DgXBUsZtfvcRnvTxn
ZVnTklbn9eLA3TqauQpYyyAUyqLx/LrjpIZFNP2ctBt6K18piXnB7FxgtuTI6udRoDlLJhuv6NoU
J5sFDdbxm/fxb2AUW2b9r04z/QaErV2gtTZOaGUhsZxCweBzgZ/mWIT8NZ46QauPpzbIFJCtAwYb
38tChHR5fkGtBKghVRc5osr6g/jFSOUe/vaNjz2WxqYbhMzIjj2tdeiQ0rYFFopwZNErAFZBOw8x
9tMAQAJtmDM0Aw/ymYU05Sdaz2FQOBxU/FSF+lCjvLk6UxsodCoja8TBkm7AnMKiNSp1m1eWoXOT
RU374Q6pMYFwtsaDCbO+7iNDCZ44aIH3RSOB4tjK8cqMSbfOjxtsEmOfUR3Fg/AH8SaWpa8HO2kF
vZExFDbUGL0ggSOcq24dMiyZJEfChShnXs8/kkVck4h6mPjbhQpsBRsqpfzPz4WFwRb7ud+TGYsu
7Yd5tN4eSavV4xLj/4EZfxgYSJ+NE0PA8dCox1eIu/IplrXFDsT84KXsnyNobO1H4jfX3U8RTJAM
gyUFeOjXnuNPesXRqL2RIKxtbCOSQtj+MQ9jK5ZTjjjZ4ZZW9895HK/4uw08YZRP7IS3NFexxkvb
TemcXmSgh9ZUMO7+oz+NINgGQnEUFwSlzxLf1tqC5toNPzZXYMWtmnjAXxBzsgA2IjQeaC0icrWQ
s7JmsNoShZUC0Vwm6UPlb6/+5P9EDDSdWbghLSHgeThiMWflCvrh23a6n2Z6HucF7MFWfDNJSklY
PgNXS7wg1YXtCJnyDHt/ztvpoKKcP6zD3sHchgp+Vl0xts7CAu2Vv9fGgcOTMsPTA0UhGgEqNDje
fQI1Vnrcd7Hk5jVC9pCMonVhgqsZftb0vqZe6zxUZKB0eYQA3KagQa1VebCO66ArBcbUYqlIFfnk
YKGBJXKIccO7pdho0yD267HgS7GcDm5P7Wc+NS96oCnH+ncEaQxLIaxNEpEgv/EbwRIA4By58ooN
QK/3g6HxqYNlFDcHLUDtLEOPWFZIN1+0zfYbNsOancAZFPFi4KfNX5G60AdVDWhqk7mboYhOQOQW
+iIIn45hkYPJ4jZRzOBUhWV5gpxzrarFTSNAybMaSrxoKxk4jgIM8IdwC5D+ElLkm/fVCJV9DHHc
hVrJrRv0iQyAlfku8J3FDBgqPXGmOAD32EySId8AHHqoJvxrTXQKx1iFT3JR2Alhzz+LI1OGc/an
pjDXjZEsj6GiNlnZIIM84QnFEjX+QsGWxJI4ypsBLeIsrRqO/kZYoJbJR2rMTbR4HDzVMG2LMCGR
0VtAJQE20oWTmAoAGVUIAh8l4wCkUlHDTHMO0xHRKQtjQMMOo+H6QqnII11Ud4naQpAUpqWBq1aq
StxemV4KI4Kg4X7N5UgmeuCZYkn6EPFRaTAdBW6bYKEOLyWpJPuX3CfR397YPAXJjwy1xIn4xwHB
zZfET00dO/ALrHihEbsXouf+N4NmYNHTBfiKa1d/vhdT+uTFxYZnOM/kpKwrdTm3mWEwHBIumg5J
Kziv85UmEYvmBSr2+TPEfWamWmVnzmbV1yt30J5C3wix5JIayBRxa9Niwst8T8rP9q2+bLxzQdD9
3bPkV5Ib97uZIg0Y9wxbGRFAt+lG7hWfDWnzh5D/592St1gvyhUaCbcDUYEe4iv60IU5kjwtff4U
PcjS0T6LC8IggXIOcdehWzEiJABhpYP424/emzF+A0/WET1cwOVwFOkyw0/T3P4hYb66UyvfAxIV
J8GjgwGm37qJXkDsrAfLril8E9k4ewQROexRj3mBx3orQyKsmhXPpIkL//FwtCdklO6cIkHYjpOC
zydKUoGjKiUt5FNfOVdHqnfsy4KJwts4Mk6hR+WxXaRZVSve+ljN+ksiuT4sQ6AMNOCSdDWHfBiK
e4cJ9D4YIrZwNwbbY5sawDs/YzZaot5PboMB0usug3Molq3g60Bfhcz6mLUnOHaRvFvogcKxIllz
ltVmKX/Y3ggrGd27vYUHG3rpu52mLZXbZh9dGz6e7SmDAPe/y0Z+vsqqw7kZnK/FtQqSlUA6ATqq
QsItDrcGRHbtV44k1KTi1O/mtqsS4rqta8q3O+SprZn1NDpV7zfvSqiRz0CUNFfjquCAJBriRSe8
RIGb19a9Ty2vTIDdv3fc+K2QeIes36bLsQIhTrntyow0wbhb8xva36cZOYh8Ph0bj5cEWm0B8v7r
5K/GXBrj1hFD/1TGO4kpx1Aulzzv2aPeHAnUJ4rGdiRfuNdtk0i+B2qzI7B+uZw8hpCz1c1gPe+d
j2hDgczwdduJVNaVXFlpoOGf/y1uV8dusHKFSgimAw536jy6gKqJrF0XtsjAYrOtbmCUsGrvZ9Wz
/fIYzuoL9vt+44ju6LT24m9K2Vz90VtsErC0327oR4b07jgG5l+udE4SxW3uD/de/Vx9g2ocmlaZ
DLIgMzU5biEe+NMqZmT8a45HbeXMJcB4lMmk4OK9z6LnEi5vXe60MeX1hnz6PVey4gc/0VMIA1a3
ktjZFor6AIgXr9z+iZbmziSI801r8ogvxGflLR2tBInXItL/DWtoSTMqdSXLI1DZaL2Kazp8ubtr
muP3pmNVRfaBK7Y9prGmYKxTEKI8ZtZ1ak7uPT1F6rVHTgyYHTkFzsDOyIPxzZL9pEqSg5rYK/Tv
LpYCk8AszQpCgFWtLfZg3scd7CaU137lHWqS4AWKIqTuBg6uE2ASz1W8JuyFIe8VydKGNEy/esEJ
AqK+ep0IM2yzJw81sbqezS1umWrQJ5Brqeq7Bg1bhcLWk98XQ1GSGGTsu3c1/P7Zhp99LH8lMYMe
LPfSP7Uq1SYrRRCrG7nj7iqu0zBFHrsgBXXSKu9HmW4alaKZXDr8q9+Th/TcO2unZX44ouIjtl9t
m6gmiVwrpIOPXG4izlXkG9+Hj4MecDPaNZ1H2t3UmvZCFrnuXxnoQUwrxjLwUh/MPyPhlTJLq6De
KJX7BF0cyuJLglAn3F5Dxm9J5zFx5A0OJBPaZhPkGpaXpNbuR547rCKs2x0ZuNnFqueyqlYU14/1
AaEQ28CdrOyQerPu+Y+0tn8INa8BxrfibWJUJy7vpdLvVI3VsTqcEnsf8OgwYv4Tgp/EH+SDKEJn
oYBq05HXfct+HEjYXC0kSkHtzSgWZ0OO3TBJyjwKfqBYs2dNWO1MrAtO99lch4khMejKdk5tDGNB
1Td5s/WyDZCCUrD480Jb4tKUHHiFD6BPkaPONnLmVVNrgJ2AFg8SR5nRfDHfUc44NBkn1HGSi/Vj
3/lOwUU5SZSWJxXUWLID3e4jxNtzeytqY+4C1HPp1lR3BHQumzew+O7kIY3xWovjwHovRESMIclx
7mGWH5snPBoM7os+Y50eSUXA63lv3BaMc3lVR/QvdXN5Fy1UhkAuQ3cohgm5wvTEYk3ypCw6a7Dm
lwPb6sok2dBeOdjVOiZok5aSjc1U+BWxaTkP6z4c7VnPHt1G+EkXyabPCYx5VM0GwKCkABAz357H
eSThZV364AmTbYHgxLjb9TuawHeFrTaRJ5gcYW97Aj/tyJtC8DEvDslRdhwv0djb55RDpgQjK79Y
ZJw1Zn3K2QhsnYOrYKAo7VOZQn0snPUJAI07qliDUz+FzesTbNUXdckvRCeG1/FDUrzEw1RUm255
QE2Dg2Cm/VIkS5yDj9zrVhbzKZd5JdIYgwcAMxkdWLzsSoni8iJ3DSpZFnv8AdQra+JV4rU3e8XO
dln2LLbIGBqoNmI8rveS/ZOVj6RLurDPTQa5jTnNiFFBT3vwmOm64WlhPTT/HbpR/Y/rr3MJi2JQ
D8iXt4g+E97SF58MxTXBlJtq2wuVn180k7VT0VddKmv3vI8bzNWx7hm0fU3KfNfA9JN3mKC8dUsX
cDioUeqq5Cp8SbaGQavO3vU1LJhcR1j5CxmSp2i/tJ/uRG7el4yXqIQPf2P9faxGV8DCkoo3EtGW
iBN7sdSbvIsFBgpJ2VqEpb2MWGNzyIeaNx+Ev7pN4ea2APcZmjioqCFz9zby1oCtYSnFzjV3jnPH
T78WXxK3xsz70GP8W/RUBRfkeaUyicbP4j3awJvUTAPuzsrVpp+l+xqeyKN491lpwuUZHCL6LFvw
YTNJ1X7cM1r0bvOZcfbiVCp5HZrslIuOTF197YZa/bor+O9kISGJf3939oGk7D7amcciosOl4lgP
Ll9GzWjlPCWdnYmmLMrZgBSnbXMWOy4/S5AfVtmJwST8qzcojJqjhJJsfHEkWfE9WBodIOf5hK8m
U6PY741Fe9mif2y8tG3IGcf9FsZn6BvU8ydZcHJFwoKRdQ10QwIYIb8FU7IqGtIBZQenWRyKimUg
YwaMIhUoWNdzMo7a1rF7T2SpUw3BUF3iBpj0MlsTsSRasmdSp2zF6hXvVkG5SpUm7Sw4cnDty6Cv
9Z2TQSSiwl2Pv2GQ5bfnOMR7BNhiroSBkEAMxb+UP8vJhFFEwzaxHR9NkSkOcS7+XFqTH0Lj10Mj
MzDZfrZ2xwIIzucQ7dGco5ha6ljQl/EZ2Wb24ew4OEnLg7xPL1ONr6h4j9PZThqXpSg+Tb3Kqeop
9AvZhC9ZJOTibKCpVKAJaWeLVz/0UlewnSOwl0Ol+jNhxj8F8Q/2BYqndW3q4OxuC7s3sI1TDQ3G
tUykLM38cfZADQZ5y9L79n1v1NQfhu728Q23QPMJXbU4lfsB71+jVbvsrWwJkxUFHfd4mzIUhmpC
1eoCArXBWThv4DhQJLNqzob8B6q1yHnI0e0NAYCPsQI57W5h/n1jPBZsatq1KdSoPyD/nXJZPZQ6
mWD+j8DMUUOCdpi1KJ3AsZKiPYl9I9BHZ9fgHbgPmLTH+k1k+i143IJZqIbI1vTwSJxF4euYf9sX
amddFdszr7DuxAGm4p+6eOb3AGH8v1ZBiocbr2wDZwkao/uP2yEtdMKlvea/cRrLiCo6tVtIkXX9
eo690k7griFx/YAtFlFtrV9CWm3pkPnwJtN/A7gJZce2lPQXw+H/rYsY5aFPD0qDSMoV5KmU0bVo
xTgejIupszlGxuKbu+gMineHtQxN+4xGcC0mJCF9cL7QFqR/jJVk7bYwxIZDw/9DtVNembdVIBRa
OKPnLAmdnvHURwjmD1GOw1tFsbpZEC/9ZHa/4uvhIcyN/kpqppN69VnyDyw84Q74opvbygzU3qNe
2HX4Z7hdpDSdgOxx2AQW1RJUCmkIH3aj8PS87R5JYHvdm5Li6oJ5feuolYBUr5iT+38pmXYraZIN
nhE1Kaf6qhGsmSPqrzB/XSNeQL1l1v+2n7RAX3XN5FbLUCQL/KDx30R9I9vEtZRLhBokjPPnSUXP
N02L7lWfK7LyItcN7cytlT/diTMMr1GKBwmnJ4zEEJXnSviH//ZYWC5W1oEGlzBP5fx8ueaA8foJ
hXjl3lnH+BHSAymR2k3EZ6ZR4icbUpKCd3TatYsFk/STDUvWpwjltKF+i7PpF7QxVnHd96pbapw7
lBvCAeipSrmttC/a3MuklPPUViC0JpolqhEdiKV3vGnpWxePQwVAdUF+kuumrO7dOJ+fqK/KIikV
cchdi2FsVb4C4dx3EjxXOknFKiBNdFlDJ+CS3+UTf1mxSsaQQ11iiA9pJDIL2d3Mptwpe+QdjTlo
4n0mhS6P79uP9fOc12DUYQX/ghra2pOXUBW1nbDn8P9SgCGqqZw5jhZumCHAarqFXLxnyUcp1CCk
jP2S6Ib+pEbovMizsxOq9NE2e+ihomXovHn8ZdpJ+F7jgZahJRdy/8ouptQR6pQC7+wHvF+/VG0B
/W6yKAo1fbYPT9XY3L5QMgheBwEEG6Kz+mqlaPuVeMKK+Gb8+so694zo1cjGgn0eLCJM11cm+/lA
hVNf/dfxNIalScnuy+h+3P5qGruudzYbt4K4M5ku7t3/pRIV5FYYBFQbE89Wq3Hv1Jf74u/MOCLC
CCsn6uKwVTY8eUQJIJK8SO2msB4f6t72LPwT8MEYZklQubfgJTDrmW8X1AWfesnvFrTfm25+DnKf
sAom+ZOU9xZMqF+5sevoCehR1MSIYVYG9TwwaeEuIZo9Bs9Nr//nP9S0g6M7D/YQE2EiVaMx6jeg
7mp63vPtTLr56NpbF3Ge5kWwEagwEjOzHLFuAihBOLuMK5t1i8T3VDcBlr5qziVw/6ATzYp8A1iG
yEMySKeUCQLLdsFK8SpYENz6ocAJBzQ+zkexBu4wzZXv0wYVunhuXK4M1nq6i4iNXledg9ycvwMP
65v0TQBKPfmcP2WefHxurulSUqs5UHpLhYU4ypKK70DsWsDYd4tx5D1j38pooNsCTd73DGyYuJDc
ADYG0KP3RV+zpqCwlKsQPg7IiCkIHJQEu9FDJLYHV2PIZ+ct3zSR8q/rzbGNCa94JzBtD8A2MWi8
0HdIsMqRHghVcYQJ4n/ZwzT+oOK+lYJZ+bDyEQ/9EGvkrHgPkwX82D52/SNTSrn8Q2uYnAOmnOXE
Q3bJkrFAD5MdB8wldpwfgjykbw+z4iOcYfY7HUicuxK4SH1aj7c6nFSAkZ9fxzvhLv+CabxHYvAs
FdLTEvUHGJDxpEiCOykXe1ckKVJQFGBLy/alzjK4J7M3FYPnFMNf28h5u07RQ0BOWhiBdOdgMDR/
7K3z71pXOcM62f4AUCmeaACeGr4UK+wQOQY0hx+pC88iYy9qybBKzGBtTMHH1j5Lx64PsA2EaAL+
TU9XbOAvPSQ/RDX4lkuay+UXCdkcU0n/RAPGpUAuExaoRH6QXV/illLvWpqNtmT3kHnADrY2oEgK
mk9VCUwgGV3R8rU43KmpaQIq/D7LXOJONB4a7653+28B9yPEly4zNelXTFIXNZE2afO05XYtOrng
r3Lb11atKRD52efiUR3zbFzw/Pv9t2w0CDQJqDfov3UeHCBGUzmobNt8LXeNU0Opm/3BBsAicczm
XHQzNwF9fHLBww+Ll29nzfOltK3JczUNTW7VKcbysaRliAKwwskRBBowG9/tqLfRDN2swXzFaXIi
OyleS9RNCEuwMnYta3rlvbOaJ4dx9nEuU4VCpQcHyfHlth+Ncg+v1/zLT5rdqX+wGWp9rW3eQ9gS
qLh4hddSh7bTDcVb3zXGRjELGnFEIBnhw7yVpkTM7BV3CYMttLSInTMy24nJZvyohOHzh9ovv4Kv
tW12/t4e30r6/blE/JPofGS902AZsusScvWL2YkIdQ68nwmgdE/Ra9t9Cd7CfEdjqY1S7R5uGqjx
WMbeaVn5FHpiVvLb+1e0tFzJD0snqbIDciK0o7udRPKjKORJ6+mCKTm6LX+JBoC+Q47wRvfLmE86
YgUj99Hpus4ymOf5WXioN/nXgQNEnIA5e5HpKwvZRKVDcPzcemVmq8E16A1d40riIRmzxxqq6pVS
Oy1HeeS3eR4JcGh8VPXrT85J3C8PV6ftm0EHTFQ8VMgmeGnP9P+h8999/L8g9+Z8rsQBFUQX1e9T
nSANX6Bd1m9YA12201uAZ+zlsQpTa4MmmHslyPWVoWYmjsqfmYFg7V0wMH1zqzCmJUkz1CfS1FgV
zyrQma4Nr6tLovjaSUR+UYBqWLfYu+uj8+AE/r0mii4a/t3ai428sJD25z7J9V4eCBkOZvISZ5Cb
68jfOJ9TGp4mquRLzhqMtfhvfrL0o87tSfEpmb7tEkdA39gQ1KnP3F93ZatmV0lrg5KGrQp5ysEr
Qbz7zhWiah4MqDNZPTKfsLqxcj4WMNebWMDKoqCda6HFc+PxPz3kWaQjHDhec8jSh0zlH4ROtFCs
k2MBBa047iL9VsYKSfB3GvuUW2ghCLDPUvQ5M/7uFM+J2lPY+d6EnCbseGnaTG4LEIfuMwcrmHVS
19zfOluwVM66NiF+beFBdlsWq4qhtFKdYC9XXVye5kkNfBC+/jBqxOpD8QnWuRfXiM+YLHOeIq0Z
/47SZ9XxH7jPLIfiDFM338FK/IL53HMTUQ9kPoMfQR7BsLdyv2oYkjmUioh8P68GlpFsLYhg/bjL
v3jhzOPvb4keuGysdFVaHMo0n5/d2DQQmBDjypRUD2F9HwDjLq/MQvi/MvraIGY/S5aWP3y7Bdy/
QBF2b9IspVsqBu9WYtxzm7M8Dw+qruUinuUrsJb4bsdzWsCCAcklmkPRkjCasPKdvfO0KoxymStv
n9jm4VuHhNg21+djXzqdbJzycdUaT6l8XmKNBdCGzA82cx3SvG0soPbL3v7/z2fnnexYO1xiovmf
X8eX+3T4/eqovxZsY0Ma4RaNoCaZchEzedg3Zq1iLMMj7OCPwIfpI/SZChj1940c1QVIukgdpKOD
8+bObVZyW9ZbcbJ9myQvfcHVEjQjQEZSABn8iZ6qa6GqIscLMsnLhdBtm2WKFXGnqklKzK+/d02A
KZVNfby7cr52UOIrYo3yRc9gHpWHCB7Qai/JnWMZjnuGBh+B1TxQWBj1dTpgMtoSuFaDJKXjOxjG
k52xT60XwpihMIVHiMcv3i+IHLmXITAgYpmDm8OPLeAithfNEoI9ovHpKbHxJSTuCmo0Yp4lDjA0
4v7xdN5X9pCG8tNHDobaskR1DDGZusmzFTidoCR64pkOGxC1eknUH/AiF589xszrYJD/M2PitJLo
de6W41KCkgoP5Ou2p+AY5nn/RaIj4DMFvS+tk0LTnJqCnXwuOW9iKX+tu1r48nldZdQIkFwqUZAq
Wpc2uW55UDgqWEHnIvQzb6lc6zdJ8StZUdqpcYPu3wUoB3d5ZRTE3/e+WNJc78ltLVgvbrFyMhvR
/efk05EQBuV80s/wbXS/ULEVAd7osFoeAmq/XdVQXrh3rmge3GPJQpgP9JA/sQ9AX+Rd9qZf1U63
r4/aFIlu7qQO86lJfJSA7tOisSxAnYKzd+ZW6lkNa9PDIeVG8fldxT5GOoRPBJwW4hXUooev2Tr4
VfumYpbk6CwmsrAazY7MetntZ1EDozB4NvSI9lCZfS+HDTaCsWIMypVZ49rg93ar89xmvgoJtMLG
35pBtiVrAGh/xZAE/Wyc1iijEGoXX6bRAAARnvdGkZh/wFA+JyWfa8XzRTlCIgrfzMj+d6mLUjfj
LNDQ7VGfaiDHlpf35ULD2WA+3rshtztZW89zpsYWu3dsmoFVM/2tqrdrA6QXGGHf/cJvTpEXSqNV
M+1gscGuM78RgrSjs4YjKxgkwrglCAO7xWLSvs5wK0t9SDd1DPVF3n8ScGAHt8BQ36xY6hgjaMKc
Bo7fXO8U/0/+qGrhHYwTcnwpeuvQ/kmOpCcGNn6lq5dp2oMupP46XoSYReKRd/L5pZMKpcQD7nvz
rQft2/IXa1NFV/59DQzvROyOeKi0NNPlkTcMNQeTd1vERf0bnubHrOLCA4YVg5RUI7cg72owSJj9
Kh/xq/wQZQVOJNbkZmc6Z9j/BTQ3nwYfaqxx1GaxCjjd9l2RL4THk4W3pLfb+JpZsihmSqn+qfFh
dp2X33q8owA7fnBSMEGCskaxiacLCTOC4415k3WVTgEssl0607c/pt0woZLgy2VkPx8EejzRSwG7
EgnlQRSFi+yrn9iuT1UPlFcBeIPy6JQblBk4cax5D6QgyuRN4ag7OMAIpogk+aFnWhBao7xNZKQG
XrrN3lUVlsJ+aMHtUE8NPKe9F5AC20CGhTwt1bWNYe/iT1elEyZk1cjm6lNpIREKjOfWci/c672H
3Y882FQSvCCpETuGg93ljjgTr9YWOEzIeHcI8b4CpUJaY5/8TLmm1NoVtK7umw6+b5ogQmfd+WMg
i4T1cwzbKeymb7ySuhwQV+5riOD1eidWREGjymt83Lpjs3xaqyGDSy5WwGwHweO+AOVbn82x8+Mn
LKFFT2zG84IEvpZJU7TBi7Jm3qbeJFQL/xFpaSQ6rHVANuBXy/juq84EhR8Dee/TxBlohy7yFiNy
ZypVkStQdZN5j3Y+KeB8wCqUDp/GAU1vn6nuzLBsjnsUAgfnfofzslLQm2FF+NYq7vMmQmYTVq1t
IhEjDFqWc8Y4PG75FOz9Eo6p4Ff/UtuuhetVMEgPKNIJUyBK6WmKXu/dbFq0dBKO1EcfMC4GbiUE
yNJMVzTcU9ZAYUPzc3vgf+zkBP5YRcnuPQOTv4j8Sz2ylzbqli+NH0lxJ5Fqg+8KekQ99iBUlk25
nZ73Kdj5CNMkS9gMB0dlTRi9dC5aUNiTqLnvdzK6btz+Y2WZfc5pfbd1iDfO2uP8FUwoUQkE15VJ
biR7jIlfUQX95mUq2tEc8qDWKC+uwj7/5q3+pLsbtnKswRsuOw+ToukT9DzNYmYsp1Lb+MnXTAGH
zjDSnYo6M2AIJeeQUAfLh/fyp4P2s7I8z8rk+kEu9utPRUaFTszsUTF2+h1ObES8lyKwQ3llKZbB
HpSt5qBHR9xzBcFzOkgfY7R/DcCr2KeQL2sErNSpQgPOxTLnTny3ialslPzuL2+5rCYM0HYsq/VZ
POFXa4AGDF+4A3EqCBxzETq8WAG6L/gotbUK6SKPtuyQF5zhTla+nz/nnPrJTxR9tBnx9JFB7j7Q
CJRC8WJQNymyNxZ0IWm6gNGkbWVtzhgBfEwiNnPUXsUwK5dz6Xp9z5CKlUzpdT/xeYAHn1MGGhrQ
Bs5cH9pGBm70bW4R9M6rdkMeWkZlSEnD5E+2DR2k9oT2rwz513L5YfUr8RBZVASFjHempkR5Icgy
F5Tcog4UqfBB6jHAkECLaJH4ZnAE8nOtlqQVTdJaaj/tb41Daa36M7tcFB0wwVXy3XENG0bIA2K0
0JCZTpQTtb77KBUCvD0so76WM+b8SnQp62TzTzyHFEk9fVMCSCyBMZNGZopfoyw7cB2vSkERCjzM
tnuPg9ta5DYC69k6/0BdaD7iS3PLeAsqXBffwwPDUJREDktWw+piHjnlLVARcTMBvkGiI/MigInp
hUHtzzzesoDUrs0wGJGO0jaH7iWz0h/y5NYrIdakiRXBb1bf65eahNoazL1HhlmzMIYvEgxfLDMm
gznpK1K15TrFylsx11Wti6Vuaht++uWd0Dt8z9KCQmK7VEiflGSFUKxHJXfmMaD41oZBXfD6ogmW
OvX4jRjlunX36F5qM06Btbtcvq/Q9O1+ZPRf/sqItqz5o1l6WycQU/k0W7/pRzwXM+nONMh6sVG6
Y8D8Qcqwyz2Izdgn26YddgwOuwHtWEQN6G+1nd2RlmBsjmfJ6gyENgxfHeM78/wnewEPrmZw5fIl
7G0T6q3NoONCOhkw8/iq7/qwnneDXNkp7KYXTQXyFLvVt5OEK/yYikpJBAghbjYKuKVED0c+sIWI
YlWQk47r8Tlte8ycuKkyXRF0H0xfgDtHtytp21R2omF85xSrrpUbyfKlXYN0opkyD1ne0XZULZQP
Wu+ZZAAVpENUMLGb2iF92nCRD4FyU3LfuBZQACkNMt44BJccku+ezKVLfsSQSssUvN3XW5xj+y5i
yPbIrswWEPgsL6Ap0cOYWg4cUBvUM9tYJMYGIxdMFa7HaB7fcsHtYM+1WfhBI9Rz1JH01Vi0qugx
JL7vuQVDYJFpx5kLhtF3tb0P89C82DnOfSFi+MC7pNrXzhdGgK32GWEZOHZYFfLGAhorb2hfJ78i
5YiuXRoIYqTn6yBGm/O1KjxblCLZ/i1CzTFGnlZSCWRCp4RjL8gNAmQzRR5agDpbc/Spg9VSmutm
I8O6u+J07wWpVuptismKiRde7oPEhX6rGn78ZvYHFS7xAfOFVB7qL25eG101Q8EBYfYq0tac5cs/
LysN+yrSv8n+67qPnD0KTtfHl0brG4hqeYgEFalB2oru1oYQdwNA/jMgESAe6tDGc5v4pi283UYI
+kkIDFdDS4KvmtdnL0FYJmrnerkKk5nK/rEgQlaKzppC4unHfmp22979DBlofuiRTN3K20zhk5Ow
mT0qajwtqrflxXDCkbBS6o5kPH4GPSy4vq6gEgzqdJmqzcm/7Lvblyg88PTzwmEGynr7FHKFhG6y
8+sProc6eQRzu+lyaUV2mPwwTkEdSU3PdCgOp6oxWr+WTJiDqnQ1/mjpb5fV8vbytuQ7z0N1OU3K
ARsLBK0cErweVaBv8f+fBtXzUDxA66j61GgZlowABkNvoawe+1c6pk2UUjO+4hprATiKkp/JXcrB
fdgYydxOFwFTXYH8NfeneEekuA/L1JGZ4i/B0db5DWeRdbUJJCBTNjU0MORe4papS966YLhzqXsZ
vmVz8SQXzO/F3jHXB1AC9BkmZk5x0lU63MXTzJyPNWrNED3USXepAieRz/gRYvipybXlnK7L/uvp
BN1/v/bYUBJWSDZqZ/fjYglfEwxgOY/N6x+yEXlGmhc+BaxWnO102TL/inbl2FljFuvwgTvzczXG
rkmiLpxES0FHRr7GBk7IIfA4PG0ju1HClVfCjEMnwURjqSe48Cq6ozfqHrsQK/eVjcgZ9fSAfauv
Yv9+lrVz+b/3e3X3DbhrHHC+6FLj6K8cUAsJ8966Pzh36GfZX3UZ3QgSwjUgRze/tsX6jCXE4bWM
3VTai8VBobOTQK1nTxfrdRtnopZ34nBuR7kUUdagXTCpA4wwf/aek9TlvcPY7UA49D3yI92sRl47
BpR6lr24r/mZ3Cu5Gq8qVwMDBPwAy/++NazjV47Px16GQVgGaafDsEkY4UyJTO//CdOzI+76xUwZ
xyYlYpNRnpzSgHu85PnXQASmVeymWfhoewkq7bIyeYsr/fJWFDIhFQGAKmmGvvPUM/yMkE46J8Z8
j8wzzfEgYqNNhd1C+0sAdSyKKmTvAiJYTezgTLRTkoqYHdtvzHor0FFQuAWdxBgbcvFyRZqkl93J
gbCllK8u2ld4Q1Nkx+EfY+6/zSSix6lGw3n4rcfPOB/u6p0x0mbdohwxFrRVxAJWj7TTe5ev6Dig
vW+zYlJYf3BczxklGN1faRy7FAZVgwLsRZ67/VOP3mNUfrzKRrDVXF44TEDV7z2BbRhEPEWnVd/T
CmE0lVFBYXp7DRnm5fFbZs4MY4owoZzL0ViLxOvYCKHJvYbA9cACTg1qg++/k9z/T4NWXA1r852I
TN45HctUrJXwZbuTgQ9sdr7hWmmIapSu/Q6+JtgH2gcbNAKwdefaEsUZ8XjdqfAfEXBXqXBetdj1
c6tfBxFnJ7kytkuz01REmuSjqmUD10HiNN5id/OiQf4yOWnaZLkXvuB431Of14SZs2JX+US3LE3Y
e4xOCd5nxja4owE/AhONNk9R2a1GFmKhDAjkZcWus+iiV2FGtfHXfrb4TNr6lWGJN6HXMNRfNOqH
U/sDDn6RpB9jGUOuTVlZt2d01/QGMIHW7kzZfXfU1PAG2wEPk+1fgR/P1MD7wPc7Wns91iFrnd9M
ybHQ507loa+GwkujVDllaldKbM3vnsHfUrFlFOyd09FcREg4n5pxi3HCeCHHO55lC2Bd3M+tNdKs
X1ax01OKUcYfe3RamBpRrTos8EISUFRJz17TOL5PnDgOPrf+qGD8zbCqIXh5OpfZzQNEbyy5uuig
wZPF1viD49xJR+NV13oq4bbaufwVNAGItEolpdsqDoZKLs4OuVEOQ3DM+WqZEH4QYGJNiPYSRC/1
W3TJvgmEAuaFEl+SLCwa1kvGI+M3YAxIyxVBGqSMmORJDEqH2JIh4YYpTOHw5xuI6dGIyp9vVtru
KLORboBVljTRunaoLJtr1ccrt4I1EX/k89V/OI0XU1KnSlonKtwLLz3aa6PhT0Uv9OEhRSLH9rgK
VdsMhwV8FCIJZRvhsw5Prpnf/D42h11bB7f2Op+vkTLHDP/3pIj/qOniVxsYv6Jo2A8YTyJ/XTNa
U/apDZ5npNDX1dJ0zPCDO0U2XyEdqjKbC6CeiU5ESh4RO4o7yeE59HrQVzZ8GWcxrooCHAn9j5Ze
grQQoylNyxkroNbkGflFJimV+HayS+Z6E1L9K2x0+bv8yXwKfCCmCL1ebPT+PAO3mRejke6emzRI
U7+hpwMkzZ6R5nSKGwNunXRgdxmtgSsPpP5YEa4Ph6LQ17YBEI9S1yVDbqJYm5pw2m7IG8uQW4NM
j7dv9DX7na+ssqh6TRlQEq9NUqRRkV+/lo7/HXN7xH/0bOXJcX5jneOHBysI7CL8c2axKM6CJKfW
hLczCoDJ/GwDdKIMb8mEO7HJDgPGM8cuIefNEqVfoMVjDrIGQWX9w5+eiRM3uWQiX1IRP6lgB/+w
1dIQY2CM15z/sREY5J0d7zWEQzT50iCLDlF0Nq9HaYMeryoVNk1tgaYZZawNtXaH7Pok7W3Wdawl
xmWFsper/hzV/LTxILIVY5aar1vJ/ja+tNgEy7LukKCkErJNp3/8Lg1Ei5KbIqlyIRztr9uwNA6O
gn1mDFknJes7UKiJjR0OEGE0Ly6+tRdxwcu5SMnLk5Tu0BGVHPzd7ZnUWaamubdnjJC803ainOTC
+p8r10V9eQjAqHmM5M6XZ9R5RfVSq7Wx5NyjepAXjz09WAsuJf2Lxqs1GPAppvFMtX0sAItHszlg
CDIxQJIs1Wbr91d9I6g72EC9JzNEQyPRSCndBjD0cdPE/YQUtxrAl4RGfDSNibDbWd+23+k2gh4N
xHTHX4YhCVhxnorQHKtO8hgWZJSB51TWkNhAOUHFDhbCxplns7lQyZFwiIHiSgL4f4XvnPlWFXhh
NmGWPVtb2MEC8D1N8pz7/ugsfnEvSAem2+0ol+qWP46iUzKcx+Kskx1X3Znu5ihMdBlDc4PaSpeZ
3kfIjg+vruCB58EgQYucrD6JzIzzu2JZweKR6ctrF9/Eat5PUymhC2KUVn/lE0r8fjk1393CskeI
qd38KDs7vmzJx0TXa8aYtozs2YUuFnk8SpA8Um9TVkgzNaCIFjQlvKoxx5H8IwUkRRA6knJIm7UN
YZXjtVIIWNctErABmD/wNsvp2Gc5c53YG7nfQCeVOVpSkeShAZEbpu4slJ9diIB8W5S46KCe1+ak
sswvhmu847adsJvHREDBTwoizOH2XOjW20hnrfWFQNJakRvACaqFR6rUHfkTnGsSOaYtOJZYAx6n
nZS2rdCWMEcQzqcTDmAyC/zTrBOlRJoPQmRGMkKFDUXuxTZ+SKK/EFHNfn522uJcrDiH91uveigR
RxN71ohV+amaXJvG3yuwRYzIPv+iDfrVUGXSuEZ1Wwivqa0WKYVvdGmu4nOZAUsmJEPyQvcMRx7p
/PHnD2TRhu0wXztJQE3WxOXDMUWrM1SpT5fK4jzr221vCfAlZXbQbhiesdqQPq3FlZ7arJqZFckA
wqtbg6fSI88Y5tojah6tdsr+0E5tlv15HhYOYcUZouJV0ERMZ3sDqyqPPF2pu3xE/cM6PXx7Hs3x
CdPD0wn0Rip5Zv3pZmWMP9FKzCT6v+LMnR+NWddT3TqzarFQj/nFpZ/34AD6ihNzgEaqODazOxWG
TNH5TLKb+zeDC+yNY8Vm/DmhQN8X3quHq1Ojj9qFBT/esHsGDzM8BrXdLhuQFz9L1CYfcbY6w9Uf
xwbqj8fSTKw6GUF03s8RLNVdf1qnbOTH+CZfVpAf9XSK+zBluabvWU8TBXGAtGIFspL+tsJfc5pJ
5du1gJ2OmBsZRajAiNkYcMpElfg0peNUxjLqaslp3c9LUN8HgsmwmmgtnvzSJhNkU71H+tg0xUm3
gcHLliPZT1EbcgNvsVHbto2XbrZx3TSxKZ7k4VULu9tC+ReciWJSJmjWuowsk9jvih2xoNFho6Pj
/pbr2VX3/DK7NM8134lUi45t5qqcvMkTYTR9dV7Av8xNXQTaIlkQTceoDfiuMVN3UxM8BFg3Jsiu
70/YSP6fJ9FgqYGfkwDQ37InOY/f8i7beHWQhFtp5R+mpppGo0E6Kb6yQjZxEMP3nMH786liLcNy
nihkixNFP3sL44JQ0Xyw/1XjsHfyZvU3eGQQQugj0OJOeOudNWcKyQesbgmQxq0wxFUrP8C6/8zJ
c3HplDhPfkR8T7Ye73O/6sH/NTarOe1kEyBOgsYDsO2dwGD+/PyrTmhSU6Dwxfil4vL2F9F8zbPu
OxgY419Dasggf5BoLiMrO375O+Dh2S35xANS9zGyY6Kf+8RmUKGA3H2xFeVrKokvBk+S2RM3j59c
D9HiDtDqoKe7KOqVu+5ujE8g0kXA+Z4VBZ6QZmOs+hUbyUuLiVtonIawS8Zj/slo0E05dIumqcwO
hIbB+2pj0ANxSFDGU15HkVw27GVRz+9DWrDrepIJobLelFCiiq72I/Ylo56fHPoYXy/tyUM5TGAx
ZfwRBHlrLTcSxn0sbGK4wDB4PEc9B5AaFCUsPB5nOsTJk5WpVidEoa2B632oxLwcpi4ZkdXX9nyt
e0oHi8EW8UrYl8MnrR5QCtRrA3v9qtr6jdHIM+C6R7I2PQeVB62jm057IIjwFkieY0AEVpLtsxI9
+72PKAbpXxHwiQDkb1FfoBeM+FQSS5nSKPT9hVcSXQpC8900N86bAVpvH9gdjHmYBt0Md5kh8PG8
e5+5CwwlS98+Hx7MUhVxLYvkFSq+Ye20LjtoA0E6VO1gZZ72eU2ZNcPj8RTYEnWVw5OnrGX724gv
WilJmBh/E+C+IFYn1lEn+9+h2r2fkwD3PmBB5h80+KXk/Y+g4JeX5IHwBcadwV+z+FXfKq1rnXEz
xqPM/fskZxylyuo/CEx0Xlp2CvocdyQKsWCFhCAaJrqlgaAk69yhlmYfFW1WWS/aMIZyoVXigcwp
BdOEiQoNclSHlSiK+UvaIixFbXsKHHCx9GWOb+XLoMciENlUhaEXLn2mXdvBhAzYThJtFSB/4bN2
FdJwJk3Bv91c3yiiObYpWVma+OBQXe6unuYHpV2ungNFXLZu2RP80cefffn5/zqxPChOx+72GG32
ouOsPyxPweBuE59riMgCN0PIMicZ3adEXlZUwt6jv/Ih++55jy9UfOMhuZ7VRE7pVKKsKRCiIOdD
laZdIkVPmIdCSGyBvfXoI5Pr43Gdv7b0nqBngIp+tnfApCOOJJMBt7XARU70tizZuxjdLeiWe2vu
KtcCtEaD0f41vh+MSR6g9MoooRRjizIVrM4j9AZkGU93mjEU8PncmXY5/ISrnhyJiV9Ky8/yfC8r
OIEWvLY+cCZM/RYVoy01dGAcXFO3X85yDhyHtaUOpS7Mb+ySKsX0VI8ZVnsZYsa8+nGWiE8uLWXC
c/5wEWAzYOTL/V47kTFU80iNZlifQknjWa4MbTcNDJxzACUNJL08rEjPzsWkjrWFPkOgxblixdJK
E+zcYIs6CPbwmhueV5PABriXV2+SM2x/BIqGefOwmKm0NbT11ni4cb0W3AufjUgjNYO3fJotINfd
2XTXEJvuMrIgU4AX9pD+DQ6V7IBd4tlHCjStUeRwdm8OflKLqagtEOLIeF8UFGNWZ0/c3sBBUgiE
L0JA18UbBse2Mk/cHXyTukzL4xTCT3SB6Z2QxuUmi7RQpNlyfZVOvsCjg24Hm08wEMJECJ12lAI3
zVTER0K/HLXfJmjTM78Qeya9cdhvnw9JFh0Ma5YhFB8RNJc+pgeoKqMFMyyZDSoRIHtmARKxuuB0
g6DJVvIryi5uD0K7Sui6ojkmR6EaM6b6HmVuCvYtixdG81oua6F2RZkKpep5igroFv1WVnnyvILu
y6E6uWP2Qn6Mi6gtNL63L+j2W+cCbQPIxIsRigAGxK+1ozvd64BWjCUmYwAkv3ZaUEOo02WEyXwf
lucfLydMfLZHiRQzRi2Uce26vZ+fz8dpO5eL0clwM9EjoE09rJYoNVyQlEnlb55gIOcJ6HTbJU+A
xthzZfIQlP+OwYdYeaic5Ap7UzBJ5xmmEIDO5whgt91Ubkz2sv8HBPOXlh1EgXHIr/wvEUTy3upb
IjxysYi468H5MV8V9eVO0REOpdfJqazwJmNLMgMVWqEeQ31hE8ywmTSjDR6DsxwhRvEMp67MXyym
3n4GsH2AC9qT4cq7wG02aAN6t+dLdqRhowX9/uNCkxxKEeiOkkp+WR2Oks9HkzhS/sI4KD9PJLZ1
prxNzDswMIOWltrJCQaqBhZKO3y2XP7taSpFM8Vld3/3+zru1iS2RqHLJ11hMU/hLU1kLl114W63
4XB2I6zTDoDmNNhJoIW4wWmpC0zmDpWXNCDJdso7AhZ/MUop1XoOcN1vnR04fa9RgpkWEYxLY3xf
a4bGDH6eQzRM6oYxvAFNUXPcNJ4GGieXNxx4VL8meQNk1Ip7KmDK5pOSr68dz8rayuKbRCWI9+Zv
ytlYaGwv+H+GkrsFY/9mE2jG7aZatd7mZzbKgCwP+8AuL3h9fTKInIuxnYmCbEh7AureImznNGmo
puG9qY1DLjIZtWwDfpdAjGMCilzhV6xdyZSFALjE8DdC444ryMjaZ0TSDuN2tHI+7Ns50Wtx0WP2
6J2/QTcVZk8AUVwZEPdFcH24VrItEbTMZRnn9JOm5HgDN6A/0PYwAlaPH//GI0+GctRfAEtodSYw
Vq9Ga6z2qly5PH4rbK8CEhmLDlg1yq+ao+MulBq0SWkYe9KTZivEODvDrYGInmNElQvRamluPieT
rI6z1REog+jhCVOGBncnWqq8i9NrtwaDPA5Qb1W9XIxTJV5SwyRdYe/+uR42zELFW6oP7Yo5THWT
18Ss//nkT8F5pIdwcZG2UEqS6smUMD8zQUOhIqXbEPbDSC8r85MTnSiPpkKv2XHexmFL0wFCYXfZ
Ar3iVTvC2WmOEyuG8+aNYiaWPp4DJZqpiXcAnu6Wxm7px0MdJZPXs77wKkubIxeCqFeCerESErqI
xf+tKYuA5c7DfnnwzlgZgxoIBEPfotHWFSvCByKTtsYk7v28x+FLsqNe1WQkGAYz/rArDe7WClGz
hpm3foVhjHDrwQDX1vayfzf9UH/ugXbJOfiguMzjA/FCOYYjQzpaT3raXjpWT+sSMczv9jiLXHrO
NYTgDks/DQ7wYigjfX7YfxB8uv1bHOoYCB2n1FIj4gNAREj4bCpnmYBfamAR15mEs3Sb1+tPqiy6
fgrQqOJvngWM+UZHEOrEcHKakdiKLcvT6oa3Mjm1asEKuM5wyoLGzoONCJMhk3JRzDBqUDR12fe6
/V8H29S5kfy38mMOFVabETwIzeJWmnrM/DT3PbXZo9ZPyeyJdaPjEWgwYKNQPaoVxgWLVZcAbtV4
53DzWTtn6I36+IXmCwaiEk+E5p5gVnHAX7Gt15EWgCOvaP9VAimZ3mIkzzNIFxC1acY5zwdyQ4Y+
ZRbg1ofU4W3KnZ6G30tBwhCJjgewXdMTfR46bSep5adTW9sBH0JmgA0gsxkXWX5ZdnD4MO0Np9BY
UyRbsEqeD2J4H3eDpEkY9JHgnBa4CrjZUHUVUAU48qOmpJK/vblUfJomAmjIYsnon6b+MP9TlMxQ
LIvYqzmZwp3o7xjSSGA6V6JnwfosllwxGWXs0vaEnvUEskeTCg2VUiLbgWTZW4JjIKTLQn2ifJIL
qTZimh3aQV1lkLoAmS/IDFYxhlSrVygtFC4NLlRfrvFooK0oon3tqyCmFT2kwH1z3QOiJPrvaafR
bYU7YqKHHDLXCsushHR1CtgPu363dk/FLe1p1gl4P5wxKSGr5oYFgqgL+yhWYl2fGNaYFehFeh0C
5J4BU2zubLDyKC/rsExg+jZEvjGqhPeDDcKOjKb+PyGahqPQWzyTRlHjo1TVb3SzCvozmfjtWBbA
9wpBE6sQIJNcA5bqfMWo/vjzmiOaMDztxbuQpfyiRQ5pju/6Kcdz1YPf6eO7YyPLtIgFlx3hqjzw
RDQYO9DLzda/zVPDsa08aMjI/DAd9CFY68RhBXVCmKeUR9hq8aF4vIiD0oVTmcHOieuQ3sOesggv
+dByL3TubPJfHwlqelziRPM15LK+an50obqGlo9UsnGuYuXFBR8AJFJYuFrb1g0tC2IMArSrZgrX
OqNN75Oy+GB0Pv6nGsQRSNPVslC+xqInbHRHgQkKFETE7sgP3GbMPueGpog96g/fDHPsf4AL6bbD
0fF3F6tv0Mkb/rdG/A30V4S8OAQuo/IwaPinPqrFpzS5jTMGnioyACDTFEm4y1eqEHFDTQhSUO+k
m9oRNsh4uhbX7DyEnG6r0C3kcymo6tgzvEqwUMBGrtBhKAudNColRvQjXl+O+wPR6G4M7PD65kch
ye4TVTpbOmhATscEskR2WGmfkmqAOgMMth9lsw5g5eHvI6jFYUpqu0HPtLSae94PX+LgF1hsIkA3
Q+Gb/4XZXxXKoZ+AKLFkbdGrdIR8KfIrGe6+1ZiFmWSj6FjvKei36dX/Fr9jI3oyKUaJZOMH154p
INk/S0WBcAxCn3aNpbHK3vLN1YH7bnqf/BdJrDCPm/9Cv+ILuhtqVvkr35xumt7OTn4Yn5mBhNYk
02KPL+QaQb363HEqq58rJ/x8xrCTibkR9NhwgldpVnBQFxuK66Ullpj2ikg8T3nAblPyTrR0B0UG
do7fwZqx4H/qNPll0QXd/wkO4WmVHqtwZN5NRHsabPaqahEkiRB0CD3efP5gEy2N40+AyVJp2yeI
mBALmiExj4qkxxSTyb2RgPvhwQY3J0sRD8SK23Frj9PqpgveIjbn0TYx1BHh1OOuafTB6JcQUDI3
5qCY7S3BLHImcE4dxWhMDv1W8OIZmXohMoDUKy9KH+KqsvI5DkQymq4c11r1JReuqCBiK1g1D2lj
LnZvSADj++8HWElBaXU0KoO9LFdAOrmvRzVTxPeSuLXB3JcHO+S0F7QQXNL4DIu3Z2I2kR1yFmcv
8S/KVsUJt9xmAQm1fcm+0+g+Xzw7ygUjnbrBKjk0frhwdd0OEdjX1HGjRc8WYg3UH1L+axAhPXZt
ScN+Tztl4JMiVgB35Req6CyZlmapHt7B8U1b/R7YaQnrhMlXfq52+o3mtdf/N5GIfkcuL/R8GVmQ
/1Ao/uyaRhhIGAQTxA1KYiUHV2IC5EsCFrGDA905gzGlmidIESQlcV/ogQQ6cVE3ywIYwQlJyN9H
w6RutjdIGDOkpUlEfwm0HMLlcefgQMjYy1YKIkEWMeF/N+FHJ4fjcJbNk7O7aU4lniT96BewfWNQ
rv3Y7MyQbFvtuSubJJRkncFu7+Vs45G1euJUUA7yHuF8WpVbhkNNQ4Q2uj2SFqRNW+X9KZPgPV8C
WDbcOUJDGtYk9OCSuPUK9x1/aU3AnwATHzczawAca+kY7n7SPSu5uH2kR0jAx0KPGrnDSdrHw7Q+
MLCEAHhKW6n80520e+ZT6yKGlBF0Kx7DYn832CPv4zvThKqkWlVVphoTDlNYjk0RRUli37KCJJi2
tiIjiklXDpZR4UxncaC3UF/gKhpmsZB0U3m0+UuekSNEGKR+7GcMW47B26bnPkqrk2QK46gdQZ+W
iiBvdxwtWL1d0Ziom4KR998rL26kEdrhDm+DgHZLPIbvJavTweVvNdiGxOw7kdPOPPjOJ20iIxLj
3gpyMIH9xxxKxpAyZxm086f5N/9Iwf0nwozpgaWyfwz2naR//Okn45cOrY/PRXhZtYu7xt6VoYQH
YgQdtUljpUWV08WAaeg4ibujc+eT9L+K7jShtlrAyV5ZmnGHCW15HnK12a16Lygexvj+YCLQB8Qb
3JL0wEET8AOG8b5SrGz9Kr+iv03ZzIjAzJvJCjC4ZeNG76PwA/Kb8Bwf7BxcJLYnSwY23Wk7i81Z
FDuJ5dWqKZJMWyvw4ek/Acpu9fyHC2l7qgD3rIqYrHFYp17Uk2ktjwXxltonvWG7KZoYK16fU6vA
3al0sb8TeMWG6pgagioiJIJNaMnXvlGRH6jKsAh0lYPnGkq7rzInpZLrNCXJjNPTjjRdCXw7tovj
8OloW6I8lat2u+4qOSfQogzZmsm9q4fVYTbckI7rnA5sne9fjk0zVxXleUnEf1Ty5xUB+SKb6rOO
OMo9gC5NU5YrFA8aav8lHIVO/2sEJv09hlybHFz8V61E7WHZIZx6okoF3zSEFoiH+ernNiX0Ni49
aGeiqxbP103LeVNHsMUgYsrb7FY/RTzbNTLxyUe9AuEjdHq9ifrGNbgg1t4HqGNYKChYkY5mSuH2
cyT2YQd4IlBP1LjIrYZDAplr349G8VTQFM/D4IKDgu6kRWx/BJQf2R1Ui7XmcvKA5Ou9cM7PLs1f
kJc99Zw2zjvrTwqWpqWn/aczWRGk8XU387dYwzaXocjA75xjBpp05llC8T9lLpo58tERD6OEsGki
E0GQK+EqVUHcjk4pG15dgIwqZtaWBJdpcwh9xcbY7ZAA8dj+s9AX27Y2kdOj1C2N7JfZrIBhCGze
TQcilJvgtEUFe+oJ/8mfLkizRKyjVd1NzkB3JSFRl6Dcy0S3GcbLZV4KUZ16kCZJ+QHeva9onmgc
g3Wwdo6dIwk/kukC7OIPVdZegoUW0byegLMUkQISC0s7csOvU0GaHHdldUxqOdtkoITxXVT4k07N
BNgibk+UdmX4jecF8KyORx7/UkS0i7CoTqxirKgbUQNLC2wyzrmlAWkZGuwMTM01e7PLBrTZFzD/
x5E6ulioCwhNvQYrkIZUxyrjDqAPJ4ef4MjgbvozBju2wCJVxvOWSBxV6fok4doQxnL7nm0Tki6q
twxMr1CtTluJGmBr+iQOjJPT3oo5PPiBUJuaxbZ+pI8pILQX/JSeLdo7gKymvJV3QWKzlYpQ+GkB
/PEwWBi058kkSmrFTRsova77izDduh5j4gpGBSck9SPtTnjnlE9OlZBqS7xfduXJkB7pZwdeotkR
PsUWv3//cJHbo7UeeQAdGW3VP+wpf49NJfAGH/NKEq4PcvXbzT0AB0z42aG5ZMjgSA07AfYeU1m1
sFCo0DgENMi4yfCZoEfMF6vbtFNAI/gM7SpYsb6mWNGa03H4Vfss1mjhSbUjghGbDMo0LjYFPOKR
ur8uF6JKXWYW9CTQi8vDVc7JEyskhDx3ct7vjAlgcxh/LbSe00mRwv791iSQQ43Uo3ZYResPFxv6
ZdP1oRabkQFOopr0cvbCnL4XxegOHKcOLs3m2HGnVGtC7QvxUnK7SzPHc65PG6DsKZ1Ic9uEJzoU
J3AVqsSV/DBEOldZV9gBrp5aTTg8yeJvyAMqnIo1hj6RlDIZuwz4KIKhrSEt+LDXGUUmGOlUguBO
n6kVzByzEoAvoPsLpYEgtQZ7Lpyr02WkejBtDIGDJg4O19pxPd8G7V9k7T2h9aboLKN4pXKKq9NJ
6sllKi0ccKcULxsgNeCWte0lEKEROdMpCUjiGtGCi/2EUvPMP2kyxRUsfBf8LrlmjmQ7/iVvxbX1
sxbmz2nLZpmPzjN4y8olAVKYDkoeW4nex0xQR+zioQ18HuwpWMuw6R5bNsW6aR2uAhjFgRLd+OcG
gj8QEFS36pSOTBIZGmG94m7lnbIcluZgvQeOPiDdBs77Q8r+s0tmHqemgsjSSeZinUi7XWgWvtLL
d0n0bS9bJLMBQJBTe+BY/PLoOLT4Km+r+F2RpTb5nr4svGH0ljs3OUxuZg1cSlJtkCWi9BJ5GmD1
Fze7lG4Cr8NbnUf1aHKrqzWgDtfdNd6nIJZY4noUaPfWsb2K3hQ3hTt4Unocm0sKg/PEVM99u1DC
8dMje09Ti82sQfkM1tBWVRXQm5kH2v1jVZT4llo7Mj4pltgvcR3/eJwWaUbwZhfMPsITJEtyKblF
6VQN34rGPTLWmKeHb+WjECFBygb/FhfJWap7u6ni0EqAqredLCSLmQKyx0rewK3nK0MFdo/MFIUK
OvWB5h5frcUT+GW49Rofly0DZu8rHTwXWkLZ/nzpZeRL/jRf/uio+Q8USOSl0Ymjl3MpouacnZFS
j5gQHj5ZJ4Xp4pRhx6LVrzO5vtSxL2WB8xW599fSSqxKuegqGquP54mjHa7iKbaXBU7m9CHocUiD
VyNJJdJeO919pT7+684K6aALnUz7kMyUjy5Zb1PeoXxTPIfdWfp38YB3kK/U9APKqKqLrB0ufQhr
iLwlk/7y8BZp9Fhd5zZKeknjG+ruEtvwrnl/uKDP92fijVUGHWfgbcxTmGf5m0MLT5y5l8VqyXOa
HxzO2NMK65G/zclWlXNGEOQFImaF+Cet6pFwhbqsJTkzUXAobb8PrCWL6OML/YEo9J3xL9zLC5b2
hxGG0GVYWhZpvhYbekgOptgvpz5OnU3Tu2IGC68tQ5DRuYP+RLE1LPjzECg1Tj6F75sKjib32k+G
9NSTnVdn4qhqXwfTcWPO+pzuK+/kDjM2seqH+rfdrJv2VbF8uaD1gFaKoIxrqmu2j235jv1Shvub
gFylYnk9x6M+BCRvJDWXFo7oULzxRKpJrSssZ82Jb98yBz6dA8lgspqO7qKjppmFnksSaNa+SOcL
ajqwjH9aaVhaOe0/7Ds+xW+Pwl9W20TlDYr1gh9tId7Wj6E12MJssXR1eBXQ0M6O9wOrfTtHYGcR
JsV5rkXKQgu+siskpk1CBsHGGXiEwwkY143wPwSPVmjppLUyqNr/F/Kfo3twEuRWuREA1R9v/kL+
BFfn8nXyozQt4s1wFIDQ3o48dooUu2hzwUxQyRCySYmbMTrPEFRKMOBJPcRfMMGgDX6L+f+lr7JN
Z5LfQZxQcggF/dBB6k/vsTgMwBTSvFjbOHKBRIkz2gYEdFsB7HpXgydEePR3HAGfSBKdTrYYfazE
KQZ9RqU4ZzQrGEuJjPnNffTcYmbw8iRhftjKDCQruMv1EUJvp0No7adrhQqcEOCtYdLMWElF0Tqj
YMFmWegWm3bqBuhIRxfmuXAVpdrra1jFNBKcn59VFAIOeQUN52tU3FWHIEigs6VKQRk9rNUb6wyK
meqBi2AwGt5LVz/0TPSVvBpTHUcQ2ha4PwYZkbOXw/z85pOepQUvzRW5tFgej4FJqoN4O3JLESaQ
mjkldcfVUffbwd3n1fm/THPTyC+2fRB/0Gd4CVO/uNcazO96TZPjfS6bq2p8HBHUpyqooRt0YEYv
+XOdS/smfICgL1RTamvqKxl/w79kvy4aca4FEC65JFzvJJXsLMnd1Z3SZBx05v/iuoU3r0ssn4FN
OOCOYENEreYnLB5SBPbBEUYf9cLvsHXrvviUrU1qQia9nPGpg0cRddmGutqNO715ycOPxD+sZCQ/
xFfIQTjhlW+Rob34QBneU9J2R3auDiAmcMb1JR60fQndB5b3OBEoU3joGWSmRB/Z6Zc4cN+Cb5Jb
autdzqiNw2Eb7APJxRlKh7WMDFRXzqo7YJLWSppg5aglCREn2d/nHSPlbne+SMBjgT7h8gQBiTfY
uM8JCdPSbmUyL39rkNG90PCGMtQwJuf80GGhlpV3LKX+MNK6FMa8j76tZMzZuWiKodH2vi7Z94aE
meGh/qSgWkbl97ZHArFLy5vOOiTOpEf5fsJBPA8PdL/oB288KMDaT4Z44SvVzGHj0Av9J9TRKg1/
V1pJ0s39lDjMYazj+dxQjGYrwndHoUf6Z80zo5XyYCmOc8IObM1x8qYM4GBszI8IlLs6ii/e4igN
r4Aw/T3cX4EdkibKs4eDnSN3uie0PFDvbDZHRDxyTwJrcFzHtO+UGa1vvr4F8wmfR/5V6O0Uw7xA
sOzddkC6vvOfYJPnd6U+SIxBC2N5/JnknLNkpNxF8pbC9MySVFmOEP6QwhEIT6VklEBD+k1PSKen
DsOyPwB3HVPx4GpWFymzL9NiVLpYAP5L+61snaIdxGCgWC+iYklEPbX4xRMyCPRZuXqeWO50BDAS
8Kz/yRLve6iQHa3zs9XyQEFY0ZyG1LUlM5VKS84tcc2NNqdha1JBTCtn5bynR+5oFIpu0k2GRqMe
/e7764pp0lPnOc3j43TRyg5eY+p5S6I8N/wdnHUK5jgSfoTMR4xX/sE0LpEiX/Y20o2tTuotLUhl
MC73FGjkQwdy09FmMce4vUComLahVoe7qOzgp8954YmrJo3FIBfB7/SfLx/akxcvTMqEVUmo9tc0
gvF/SJPzF/wpbS0Tq2lTtSR0Rnj3AE+KMs4NUJTzKWZq7DwqfXxaTxsSWOf2psez586r52iGZPEs
lgb5LWkxOqWbxGy89Po1ES9xVxqs0cNPlTpJqDZS5qeMlVoM/6MyKJwbgXA5EPGUTq4tJXYSaoYw
1H+KMbTm4kg9cNCxG7qohoCW3CCLfkpzfQGkynZbPivO7XPxvQXP0wUT9U/x1z3zlQ1md7OrnsY9
K1RAXKc3ZpSi7ffHkp01pdXfPxqTc/z8q3jdyUJ8ygmEag2siSYKfU3yNgW31ztC9ljjMiOByWOA
viJ/97Lac7XWi8SwKMkvXHNnzMpqLutr3fwpJl7q3n6NDQa0kZONZtD6NJGrniMEudOhuYthfogI
R/d/L7b1kXaY01n/UJtMRe0V/wcuEj9mdFQdJhBQrV/iXaFcm6RANBzhjSb5JCKNNWiwxDUR7vTT
ypYL64RZn+iHd82PWmmvzVDxFL+V+8CT2Bu9yw1uk67aYN6bWv+gTT+a9HseOckqUXLAKtpnrjQd
ykFoAeQ20TbGsk6RbLUd0QkEUGMZIvYn8vdm0Kq0CdDKOKusnfjLUsW00sXSD5GE72gFwN7CUegE
kq0HMvfONhRZLOzxXOfP0iZxifGhMy0OtDGSnEzPWVvseIzy+QvUfSwg1y73E6NaGYBKgDXzF4kN
If6TqttaSGfEmfMpSJMuNwkLXRdT5y6z3us4bLgOrhGZ0BUXGNlyN8il4JJETl0Lonig7PTOXAAU
oWFbQVXtKr5rsIS8rmmKk/ZoYyc7/Ua+ZNkooZhRGainCqhHcTsjEc/qgP9NSasMKaw61u2CZ5pS
m3KT40eSr1jpTBUJiiaimsQRobrVVW8HoNgJ2X7Tk9MYzZvCdR13ucnWGSR2PEQsfEYvzrHrfBVI
moZ8H5b5f40xfMrd3+D5n82ZN9yCdTcc5VkvDQnlcMGBQswTTkihuJGuGUUYf6aINHxYByvM4Q77
PpzlOOwx64vnQF2/T4MKLLkQC8/gV65kxzA4uzHdCTmzdCw3z19Uvlzw7MXkXvirz3OXHd3S9o3K
Ac8/5F9v83crcSc0fjmCoNnJtvVvNIlU50/VaBRjJcBEINpR4BLQqFvo6yX7ZHhwM8oUlw/pJAvU
loFGQ/achE3G3oxNPG4DKrTLBFrnNcsfxow0O9QXPZOdL+IMMfLci/AXSGBVz3Hm3fNi/r4MwCUI
Vnll09nbK+W9ntl2EtUM3kWA/RSw0cXmQuTx02l9aAvcj1PByRjQBSNCnod6oTZ6JkNQrULlCtoi
OzYNFFtJYn0p5dOu3giej99Pb3lPiRmw2Gn/ZP9ahqA6vDJHmtbNYojEdLDH0BmkWdxhxL8uJxlF
H2b9q1bJ0cVqHr7/h1dzml4jFeLn7f3kHcn1EZadCMMaIkkq2SEpsGX+cBwgGhKzanwnI6TOGceZ
B8eDKYxrLOfdDtQ1Hqr6rdS+u0ZN5/mibl7+ViVhtGOd5lHS6IwfwqYI+lgXs+H8oPAX3OkAGdM3
cvgfXjGTSfiBeMkkOxZGtmsAp5pAMw1o57j/U5bXw8lrD2pBQmUNl4B3OGRiY9UnmOUGRrXsBTfr
scZgY1jSTV1GDTVA1mCQYm07QeyAJqqpXCoeYY20g1KscSj+OjjGpV9/ZFEjJ2WI+rPibNQRnliv
H/DL+LGHIZ9PJH9roTgo3vrajsBK4AChQWftqpuR+oEfr1+Bl9pqMOGY3XvJVVc2u4CGOGEH345i
6LqCDsbq1oNGe3ztOBV8jPIpCBIZpQzu9LYs8BHUIk2GJ4ycdFpLoyiEBsDUMN3qLJ30R0pXPiX5
2BdVaTb0hps/cIsCCRbrY8Kw19iI+vQwKADjhHCRZMkGuWXDH0Y7YKe6ab8+C4fpu5dHR6xVmaR2
/xBFO1UNIXzaty1+qZlGIgZYYLWReQ027jiQkSQLLZlIlBiZCTmZ38xlOrXAwDphYAgPJ8PazBcn
bL8mzEDlmIFtsZSUNkqn4IdI1aQvkBLQm0Z2YEGGcpun3w+uwuHTAIF+o21ifGTagLxNeOsknNLo
397cMp7fbRB2FZbhQYLy6uWnAUt5Y/RRswHH8Dxn8zlwo5nZ6L4IktsGRLys/NYs7+HGwVtmoQ6X
M5J3h5jAgMka3V9oAJOIHKW4ukJFQk3+gJfRq8TiDsinFmpzDIyoxQDrWYMyaGEFsKso/S7Frxq6
AvfM5tHMi+vXjWapfSMdMFdaQMOHF47GtcLUaA3Q4cMvEewONpReIzxr9sX3kR8MHSTuc0n/dSQY
UozpUqFknumTdgcU8fz943sC3ez65EufGDKVrdYnHBUlnbl/GWzXXo8naY3OSaEVqEkq+i0Q1FvE
Vq24PYUVoBEV9sA7XwODydX673PflEu1qi0SGvsndN3+Zg/AxoV8q/lQ0kXP1YmA/KPJeP3OeIp+
QEA137iWETqXSP80e27HyEZZ40XoqIs2rX2ShPD9JcZTuDcFQi+JqEuQ9PAWNrWFg9N+Pk1bhE7F
1YB2zniYhtKZhUB1j/GM0/qmdsecuNzEn6bZ19QOxGSRipfZyZU/SbgIVmbEplrNXmANgUjznc7h
rV5oHiHXPGwfBT1CSrsm+u4vH4nVQ2kfKYAocE2/q6qPWCxN10S3SorXrWeBfqYnM0TbRmLxGtpn
5KNkP2nwNr0H7IS3wS+1HmmrG2gInQ13PpZj8cUtw5QMcXeJOZliwB5+F5wnVw1WELHdiSyUXxGt
D6NvK7CxiuBvOakCrqKc2U8Oh8yns/6HWbYWVxF+k7mTwwhA/f/eqWnfYN5HV/iHKPvQDsbVmvOB
sgW9PtY1QDPStK769cqu0+oi1u6vbOCC56Li6E6e7pYPRj4qhikbTbb/Yo15e+6GjqQrllYjQbZD
HIf1UjiOTDugqzYQi2y29DMOC0TiPjw1geekvTTQdOQrAft8vjwlQ2xQs9pA1tKWnc4zTdbCzojd
5017e1YAHkYwlzWlKLkwhJKwJ6hLKqjXzZ/ByydRqhtd63FCRCYGLNRR1KmytKex43NxCyXeyB3H
mQM/41/obzFKMxiywm/qC8eiHiwdhwnqbx7AFjayOK+SD7jsShviKGZ1wrwleaqqcz0N++dppdR/
Z2RZ1cfEXBwN3QyE65iVKXsTk/IRc32aHP6oYePQ89y3HOdtuJMuo35i3koNosJdlnuZvDC+uAnV
kRREmGMlhAE913RKnWYzYJ5nauOgkkB5OVDh025eu4xsNj0SFyHtsv/4/X+n4imUWq7aZ6+6lVCM
eiCahTv48IYC2B3qtPeSHS8lSr4bPbJ8w1KIqgrfeyY8fR99JFJLG60iI1mZI+CWYJJkRhS4UDz0
+PcdvxSqrmPO0ycfEC+fkhxLx4rodE378QdWuqR9uDHiAqiS9gocc6r5pdYPGfzk8lIvDT4dH4Jn
1TVaSGE6PLBu+osvfUcITjqLfPRuXG8KsHDH2mYL9yOnKVbISx+PQo9Zhh4uITlEIuPiQd/IMcoj
tX51BiD6qsX1eerX0sQarOjQTbXMguXNKT48O0Gs6iJVp7/jD1aeIlUNJeMk7uGbyJ5DSjTBTKjz
470660Gi7wvYokFD00Tl6EgUN2abijlF1t2Z2TIzy0fzrN3AuiAKr2qwxK8I+wRyNuIz17lbYHPa
JwzboSg8qH6IKHYp2JGoSEF7AUV1iAFmjIaSV7cKdQOzBD1gl2CFOx1doJgPud6QMejToJ0YZT5v
3INb+bt/yG3BdLZxMMSJ+uXb3SipKDOWqNCnp8VE/PYKYt1F1CUVFZZ7fZPMINP6XCR0GYwJAk8q
QK2Zy5ysCss7GoJ2sQdSPWSpaMrk2BdI+pTS3if8TArEXGSRjRHksrutVoZVacN3Wdi3/ca1Yv2R
MW4UUBg6TKE+YaIoeYMbPWNNWTOl02bPi2nBllJgk6a1dkSzPDqfvvCYaKXtGFdFXVgeVt8IxGUZ
9VzgzmA3OitoiQo5y1O7UlWd6MdDH3FxYI5OC3xhDFHyg9tYFjkUhwBi0hpmBbL3IHcCPEb2rGlc
5EjY9cG/OlAFF8i0TFhmQxhaaBmM08Us5lIudORcbecKkfg1aG3Mj9G3mX7uutbB+kikH/UKE1zC
4cqmAzsr8iLrdww9/ngerRj5yriOwCzLzX0NeM2uA5LQXZYcesYqZAd9jqoZY6rbNKq8zED7Et7B
Djj0FgJXRaSVwOlGf4DbcVwKESWEbBNEZRA5LVX6MDQZUabLdeeIoVTOy0fNIZ+zVZEA13GDVp/U
9B/An24lLWmIO1oyRcHqA+mra+idfIjmjcmyLSHSuy6XPuBcpEEq6pKfAlUL46Pr5ZiH/IxWPs6P
nAIR3oTVpqXKJfoUJulPCVOwqugL5SWvu/KtkvXBMsjJ5g+wk2Sdn+gh0scEzzhDngpznVHcis15
oKUZNCU2R1wmVkmfbksa31HxEX6AfdoMQup349ciii+1HdVvbVBx+EIwBEOH+fUxQue2sC3AyD69
go6w8kQ2O/RYWaSFvshAP8SzsBjYURJTq50OWfGtercqGN7n9PP0/NxHYTVHOH+VhOpA81MTYumP
qt0ZFga317QXxCBi3MIukGltwX0sVYiyrpQlFEv8UOjhrUaLLRIqrep2wwz/63PepoFG1NRORbdD
sqqw5UjvpyX8xB0xrnYVTjiLWJ9a6WhSwN5TOQZab4KW/h5rTG6v3CUz/tP9XhTiQGLQOH2W/ymP
fhIhP51ddrJRP0iqBYppMt19fThlZLYn5H02Ng+6GYUjsL7XRgr2vvE5p0DqhK5cQkoo7kbuqVx6
BGjdkw3HbXwkiNh8FCharr8/2XMBuJLmFFAEMtWjGRjGx8SBX1DzHrEPYTh2/KSLJyGknsyq+6uB
jIWe6ZkOa3GprM7BCtDGvU2KJdngOqxNtAIp2MX7HQQTf4iIGQTuc5kE0qkKNTZA2WoixZ7lsbK/
nhoUvnkCA8c8jBxNROOzzf0N0IRs8HcH1LjPctDvGuiVf2xNHVTjRvTcYWyjdk+kW2rUT5eQ16Mx
vHJ+eLQhXutw1FBp1jj8RtMdrkl5Z5L1QL1LAT/wyV1kXzWO9pvlZaZcGCgnmTb76iFb5RiffuT3
ZJ1eovdX5JROmaF5al9zsEpvHQfVn+QXcjiREOEpwH0DpB0CO6uu+22S7H3xwXfYlCSkNz+HbCWk
EGmSEErFGt035wPpj7I1++tUThV8QDlSK4dQoDpE9idTGQV4Dbtc+dcbLCu9WqKjRbBhsEu42srY
rz88M1JyO5k5Rwe3x4Vg0gN+iqXL6wLP6NJj71ZDRx6q79BYb9VkKVuAFvOodQfVvu/+WMuk2Bm3
IwplYo8a14khTNp7gXhnarywnEHSAuZBPoX6Q4aD4/2XV/NhzyAdC8EEy/HFzLQn2Qofc1zqJuO0
3uPIJ2B+PCxOEsBWOm//8QGOD8Tp5YISI5juVaX12kdYJLhboW67vVsRT5LRfkso9+D3oVFY3F/o
+obeMdZrxWy1u4vxyixf+RKaRnAksEBhsNlWyNk8BsBnWR+twDwAYKl1D79CmqHzKnnU+oXH9hYj
aE0KhPxhZJn3KoObVeJKifLo/BhOb/AveTezwDtpZ1swgWxo/v9Z4bDCo8Egk4dFzPalnowePGAY
zEQij7SfIMYk4bBCMzNb7C48F9YsmAtMltOLGd/SO5HCYMmibR/cI7rAoCrTnWAmqXlbp1HdKhwQ
gTFddi/pzkeDMF6T1uLGiBCs+pLkl7Tx+gsKO0yt5a2puaAUOs9LomhMHlE9tIZVJBgf6AIu0+2X
w13/nu0bq4PEur+IPWkKXAtIo5g/ehsiBmMGwhdk5QrMZDt8sAvVAF/yWoHYxfp8wQLCisbR4Awg
Wz1jnGIuzPL9mrDjdMmR/iNOpd4c2LwCg5YJRLYqBF+J9uPfmRvDKwSyGzHCQfxCquN2dCDsot2l
k9RoUUV7dXIeskI0PTw5ZSB4GaA4Mdn/7AOFIhd+ba+5ihkjSbwbAKJ4Kl3lmLkNysEqiFALx7gz
9njtNIiFe+O1PmcDIcczrqeaNBnAIIuS7qx5xAgV3ASk3qWkFcqGArqrkB3Rb7x35YvawwT6zIAy
V7zU6/aWCWn4NS2Qol1td0cTFspm5HIKaQxLnLorDjO6As3z/Bk9dOgRrpAxR6vs4mD566ZATJkY
csAWK+vaVV374SbwZm6L38nLN3M5MA1+0U2Slh3E6VwNAxvNlp7EUcxxufDyC9keBfUDbB3YQCf3
549Usw/I1DbyeCVTwiH64anU3Vh2hLdik5EMzXimNufYUALdA6HpyIyUHpQNhhveWf8TMI6uQGKd
o3+iXqEGz1H+PP2TVM0VbVMF5r5QkuUsxFK0Q+U0iPUH65PW2FdYOvQycch44b42MBi9OQr/fXmS
ryJpQMa/EBiC5yAmaqaJ5NCi4B2j2xAbR/+fw25NR29ukPTcs4LcLujvA48wNNG67rpoIgOnJelG
rsZ/6j5jRd5oPaJqE1ED8OEyOaoo+CYW5NCa3zNKPKVXWnYSnQvaXU9WbEHMqJt61/irUn7nBXW1
vXAvSTP1uceyGlI9bUv6Gnizc4H2fOdIpcULLZNnlQvpBTEcRs6M/gjIBJde7/0zmLy3q3RkNeIZ
nCMrdet89Gg90lH/nAzdfXVj1jDMEPVaJEjFMhW+7N6GyhekSF/PtnbYNYbboAL3TeS70K5qCPzh
wN2/fBL5tEN73QTrfCuzikpQR3jXvJeWO0xKVtLfVlYYZN1we30Il++0fIfCrRllF2ZrAFvcOOUg
SQCWsKPgZ5EmGlm3TGsvc7VAMtvLNX2STySB3PWMYBJoB7RKp3CBbALcvGt3GW7kE1aEQ43l7Kkc
Re77H7umg++vO3c8EsI6+uJtE6nB0MDFj6vmJt+iSF7Iz266Ib+bgiOU7htb0I6Zvg30aXRwwOaC
TN7bwRsr/wwvRZcICW8RBlFDV459P/yyjMwGR0MARf9jIwtqzvUnTMnsJ9CZx2X+4wBLa41koCSp
8iKSidwRb4OJIH/yxsjloZd0JaxzYrdNkBovidqbX/ipY82t1X6Bt+GJg7NwfSH//PlzDhMtYfzf
dU6tDtIbxcOmgN5aIMNFe52HvwzioL06vrPtxamzQSiVpZiPjfTPYRacdz5VijPjStWNuv7YQMrF
btgwWnzRDcMpKc7S95BYwQX4iCnucR+lnp3vktG8iYuoJHZr2qw02nX2N9971vw/sqvVkfEEuiNX
gmXW+zyI5m9Ab+FamDhnOUkSJv6aQ6uXbwsFHLM1yezYdjVRC2y8Mcv6vUUgwVEAOTaUAZ91fsm2
K68ONy+dFEbjiZboJ4fveAFriaxIuzTZJVhgDPqHJ9m/4mV4fk/7R7J2Zy/qU1XyDUajDMaqMiHQ
qk/3e2kTzdP/wZ7wfM83D6hVNxmYklZpg5oP6Dxk+Xpvk4NDJHc5NQqw8Rfj8Ydobw==
`pragma protect end_protected
