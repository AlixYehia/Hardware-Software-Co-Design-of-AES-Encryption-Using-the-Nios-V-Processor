`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lqB/ySJv03F/1cen7V+DEd87MKtKbRywmpcMEG8Uh1ipaJvdqxR5t1I3laVYn+el
pgq8VxItS83jwo/TZFADYNlDAaLaTqDndbyb2dGI7Q7atgHGRvLcgB9mQ0e/l6Ck
hOaiAds/A+ECrxVnIPNzRaf9zKZ0o8cfjLbbFGvpu4Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15632)
1cs8vkAelH4asz2qP4NNAYhz5HixKQqQ4n0OQsKSa2j+A5uiU9ocSmzNi8ZihqcQ
LvZozW/Y+S99DSGxgJ/QuFNL3bMEKtVJpFI+zgpZWq1uWAIMQJ9nA49omY54YBss
CEfcAHR8GLepXI1SLhzxe7m3Co6Nopk7Qs1lsGMtj7Fe/Yav6dEYgqQwLqDtdLwW
+BPFUiT4GOBh+k4Vf0FjpVo6GtSBjjx3kC8UYKuCZP55+kCvNs0qBS/IKVrEKqaC
tM5z6/bWzkOF3ouKHvFo7LZ5ztY2SsPKyCSTbKT/tkX2FnvtI+vxix8C4+7PFdZz
wYoZo0MnxwwuzVXZIxEa4GcNZHdhYRHDcZKwwrSKXq64VE6sr0ndgT+SNamPUANF
rIN9OZJ3YUficXrB4HrADTgQLd6F4RmjRjky8PyBSme/ENZD8/iKZuBWKQykRcZn
ssIz4Fq9JM7+tahrnE5fMYuEEw0CdlEw3m6uNNEake1zPYcmbxxXj2ALfZNw+GO4
WKY9JdRxitrO1bqoy95S+ZNNxpmGnJXWCvSS9/PNXH6WCXrrPGjHtD8IsEnvrtbn
pfKUzAWqKKEU6lOpuL9Hpj5LHrU/pNntwHD4usRsdglAL6Z3yokuIrjffVADkalI
XjaRf6NsuV8J+a56FHq1XJO8oVo5HjQdI086s0Qf0g29r3OgmKtW6lfE+zUc2rg1
LTz/vCPt1S2UCYhoROTsgeW97ei1tlhe1PuWdElxn4xlvM+kTFZpIQvq+NKwwvfr
uu6b8fzb4JjZO6snso49mT7AUr0k+evaPNK1sJ/oNE3HYKDlU1LrjIiVGzUtGpog
voYwI8uGilI5+lQkvy+2HZLan6F+sW3OLTM66STzxb4ANF56JvdIwRZrEKUPYN7y
5ahCrmrG25ooo3mmQ2H9U7K4O7MUuuIpyvE/KBbbrNJruTzvDK2VP+0TihF2GcCW
PkfgORfkCfGJe+3ofJNZaw2jSWqcu8v6o20+KjU/LVB7G9wHVQlp9kza2EqMZQf5
YMhkyyJKygRpggMEX1/jzDzD5cmmEUMO3GLImaTIgRgF8uZ5AT6RamBVWQscHsbs
cFXoLY6sGR8DNdqWWaqCz+mAqPcc//Gt/UcEoHpGCj/QreLOz5K7MJ9FsMWnayrK
5fBKKRbGYQwdfwHEotK9ILO8yRomODruarzqxTyHopLwjhKvhIA7OXjKvGcQ2i7p
8alUa8oWO5ygCGPc3K94BUVkfOb/MT8I8J2p3lN+yTymIqlHwCGO1t15lZMYaNxo
7QTgjqlzK8nq2EnoQbLtkwhadOHfi2zDmqwrGFIQAD/1VJhUK/DOMyD/0/2TS7MD
500YTTsuBPvXYEUxr218djHmO9uNmM009Ij72LHeqYWH0XvsFTkf+iXo25kMFr3q
5QdekU4EJJJoDpXh4d9sYIfPT/8RQZm97FNZbX/AHOF5PkqbRI0Fn0wJPHhAunvw
VGrcGezTnXkv5A0uoqcc93yF7b1so0BDSXGw9hghmuzdCv076DsXP7M5lI36VTRK
39ZS87Omi0fOLL8nn6Q7/yEmGZEgMJgIzzzNKyKCdJP7ygFmVNyvqFH6OcesRf8F
ecrQIzEpFZ0rY8VLU78TEneaYHEhLZckyb+ozi+ZP7iGqe0fARAFNf/jRCpIx6gE
DVRUIXIbzkZUuftn1hEGYNR+25148Al+QQgE9uZhKiIJYTY4mKaHoFhth63OZSOA
Hct6lrO2MdEXvrHM+VDxF5kdeunPXA7VSYnIzY+Huq255sW9CL4uo0Ot09cvp+V0
A377l9kpFOXvCcoMMtw4j6l199mp4EWFGghs+czIzmFPr+emAY15sXZd5ygUdneU
LeYeIKtiwpFuAIK5Io6KRBJe4CA3dkHXihykw10krSh4chR3HdewPyTVSzCkgpZl
HknF77Epn29WOr72THUsdFmwzM0xkLSD9DEXUxb9PxtXTf7d1LIsR0BntuhLQuX3
2gBTiUr9UeB39VxILbsSkcqaOtbEjbdkgyE5C39AwTFHGyRp/MKyUynclyurCMbw
Xr72ybCHad8TIq8u/AxJsXU+nYFJtxfL4MihD4UpPIH6NLCLRZP8heo9+k4378Wy
Yp3vFTcrtSxHfdxhF9ucIa6R23YCFo9mMD8JdYHW1MBR8OZ9bVrdspdV47s3RxZA
WoORNnNBVPtmoS0xh7Cscx36qvVJsNY/ErNDIcvJut91HR+9bmfKj9PaPUTsDHnF
84sf6EI9koWblX89vsjIzMXxckXXuP3LDB/ssfesKT1yPZt4TVCPCjq8+O74aMWE
hBVWaeJXK4HRt0L7NbIvbA0Gi1SDUBi1XqX5ePi7mWZtqa5rrBlTyMigAOGaKYJC
jqLcUzloVdBLYtHTPkEBRCJktAs7r7vO758lexzn6624vJy9zFjLLrmNqwsIBW9j
AKtk6batWdmm5e6fUENcNP+YB7IlnwjhnWFgGgk9FDcFeCPB/Ztb0g7MdRbmoe8H
NkesnCmqwz3gFH4OEU9fXwnqqG6KSVjKg3Y+/iT7v0mnxLPL9W1oslkO+CJiiyLF
X6n8wezyiVtiXj3h4emIX5E9LiwhmJ+dhSDOs3cU0N30RGclgmMjyGsJF4FBfos7
4sn0NSJiWwVBMMMUEFx3eJkYhzhL7fuR18G6tT7ggIcpC39JLopn4FenJJtHbGdO
qHus8sUr5K5u2qqoORBw124xkg8/yyeZLBOpq+je4+eZYLwy9njZrH0JeubGY6G3
rVwjjrA+qC7bAmUK9efNGdvtRUlTcI0D13XuWptf11NSIlVfN2cuC1bKsLDuxV5i
qKBeZL9xYFfO757pUVoii3uGGzNPMEAUQxS+tHXatr9oTRfcPrbl7HBMfmvVgahi
CHkqBDQBXtxeE9ewmpbkpTX7qB8IT+nCUJxAsV8OmSiDJUMnIK8hLSXmOZYwpvGM
AMSLbyCn73vMvmcLHOmUCcJc+V66OD+fyefDYg1ReosWegOQcV4cj9XMkOgyVGfY
GNNH+KCIyzxF/VF5gG7Yn3vdhR13m6Y4xUavY6Ks1oaT9Ysm8tQIgSMOAVHvF7vS
GBdvu4fb/IPILiGrAuxevlTGZqanAaRzfLmB7nQJpwR710WMOuhR9oNIycTRxSz4
5gRZrxGrMg0/+IIPAoGNFj811zsq6dfIltpDy8myQliQ10E1gc8GslGp6slHCNFe
2IM8yHM17KR3YR8aEdlnoFUNO3dggD3vrna1vCy7qIP53eeTwLe2H6CA0IabMdY7
oT9LF+VvcD8baI+BiTu/NNUg1qEkQVZLPl9dsnSSLJB2DppiN3feKkO5+UI5NWkm
/jmJZxId0R59STTEjCRlOub/Zhz1JDqZjKYA64mRpZ3aUdRSP+tvIt2oYrdnxS4M
zgHgYBs5/CNHiqNVygUw9EMvonSAunSCOuvjmDJGq42gMoL5JWBgMis1/yXCS/i8
Tn8fjrpCFZ9aJlZjhkJdsjHA2f1lr3QUtnooiHm1tRze5ID2UOU5ixzm9lEShmhB
d1avmJYqMZ21pdkf0p9mOMFv2kkpGiygDyob6w0HFqxNBz+Bm127YFFSw7nbN+bT
GXTyxoxB2TzM9Hr+sC6PxiPHLmV9lSBi9tNRYO+3GuPhZ7W5GttSC9SucqBf9w2j
xVtCyRck1Z4/VvTtnUmgKvwE9LOaPO8doSM+hr8vqSAu03SXcb0mBbhHfMQ4Gm+8
q9ebVcd5XzAjstWAWbyt/K7BKXvPpUwj1og522i34CB1riBKRiG05ST1tTO5qX23
Se3DLmX2NOTdEQL9pyzcRn18wy33c87pUCpD3tbMKmnPQaVxnaYeOjaSJrDdCx33
CFgZQK2eNW4u0zW/Pxko0qV8XL5ChuGJudNFTyy7gZ6pF7MPH2THLYroZ71omukS
ZWFaSh9XjOnzz+TdIyCHa9WBBTmNwVZoKKxtodTwQL4MeZ1+TRKxYcQ86EFRjrni
MCccPwxpTogenaEFXrDuQYtws3lwyEQYymABlFTvMCbnkldQrUHpBvxWifANteSh
zNPBo9YvDNf3VloF062zPAoo7v785SSg/EgqNhyOvJHF1QNeQ4ry6+6BYd5s6391
DYgeVK7KK0fHw8TJZHO5fhxeROABAZNigv6zRWy3JcZIMMoJ8b34xogpp4h8EjQv
XYN3p2+HQzlDWDTdRcET2vtK6i1o2qWurJTC2AxQRQ7b3pQMv8bDuG/70uIlFy74
VLR9NUhhva5onGisdL6tNE5/6nWW/t5vEkWLAIOZ6q3gnDs5g+wkLshgl4qZjzYg
zqVNtRiLxqWyyFsEBmAwptd5NtFL84RAM43nO/PlJhGg78XUc95kOeVqAyvP7OfW
g2HyZ77SprXsybl5lblOSn6ySYLf48p1vcGSwiVOS5fa8niRQzBL61Je/aMfL7xH
GwjbfkhbCDDWkg1aEJsCACkMEQhabw1nDyYaRmbEbDd7uvD9gUPdxYregVtsvh+b
+OwnZu+Qo1536uJ/+iACs/luP9SZP081m3cJGHmExfj8WvC44TMBWPmCRF0pCmP5
BVYchMSMOShOvlXHXjYRZui/ppAxnotsE9B0Vy4dItJIK/vnnY9M8O+0F/aeKfQR
FI/kN6T0CgQeBSSRO6032G941ZtJmCalKzCzQhSr2KKVUjbXK7rJHLMV0Epyq++P
dP4f5OgL+RXO5X5N2rTtk2yHKZkBq5sDBAnE0RN1E0gPjZ8Z3U0cA5NbK5UiMGiq
Rh4AoZne1WjW9iNCj/RnGT2v/SbCxlgfbeE/oXHPLzft6MO6vJLq/ErwIcRSP6d7
+wGPQRGjuQDtndV0CSGY+XnYKJNOEcLdPuNC4brGWdiRrYLgYxrJBGMAgt49qF7O
UEBWKJnGR+4kM/b7lsdo7/MNPlKbmohywTQBBRl/x2I7tMEBq4yM9t6qgSSTkhfx
PEEzveIuwJVASIF0APg91h0zQi4va13gWdG6AVPdNXvOLygi3NjgSXFt+0RokQje
HGTq3Lrv4itXsncKKF2z+J41AWHcV+iv26qjLK6aLkquPbVuuf0QsXp51XxH/Bkr
yadgtUg8KZhsyGYrBkdW1/W2h2CeYZTkfOQrmBYsH8jrNwhv2EeKqgtWfhUhRPuq
3QYOjbtILdtHzYkAwGwlTdiU2DCXprPTLDUVFQ8qpoKenbYNdz9Jfbx/sa8XvDwm
FMcPmy2d98pC7opTNMeNf02hXK41PZhjrYifEZBOX4lSCQeTnil8J+vTtwvHdKnO
CLqp1CJfJM1163vRCpIe1/c4+s9y7ibPvSj6RcEhWuQuiPZzzUSzEf/6VMjis1sz
v77GXFU7r77wNM5Lk39H0IjuU8BQ557STxN0LmOc/1dWxNVRssUkiNGIhoCvG+Re
ZXSOYg76KYkfSrCT3FIlDSRUOKhA5AxO8LpJJd4cuSLruVKs+4bG+A95R4RJkz8I
LiVafcUQ5iM4dnodPKcTBSB61SAzBWza+l2t2d6lVuPKJWAuU5Dt2jbohrOdsTdx
nS4orqkLS58zIP0Gj4F0AaQdFmHllhAeZbHgF/hFA/nr9/RLPIlCidL2bX4mBdtg
3mwpqdYIZmSFkyZtHJtR67J1mYv7qPhNT659NVYzLtEG9rammT+HHpZOAtkQEaMJ
RK2n8wId8S+Bo5SCJajKZXxdiZrFk6SxJ7DQGFctXou7kINuLE/AuHTHgkyQ1kLH
Po5E+UDS1VNhjgrbf7MfMU/I+kNN4WDF5irDwUnapU9vS/OhXoqeODIukPsa3M7E
QnU8IBFm9XAz2E8YZvHFtn6YCPkD7UIDZ0kUGSbGvdFJtAUKf9XM6BdEQAOw/CaC
mzmZ2sxA8Y9/2BG3wjHcwF99E9xrfSn4CWf57Er+b4FKWS54gLGsgrxf+4CAzOYi
R3bN5Iqxjy6g/QkGPoQ2I30Y732Auy+YgdPKjxGCEUmfIzbev8jaDi6L7Jg9OlES
bzp+TjZCYq4ZfarnHenBGNdIji2LqcnCLSBlZf9/qIyoYyPDRYenznrCStyXrmAx
wNg0gGyjFG5Sg07IsE2uLDipFAekIJUrnJcTc91F0fMc12okrnR0c0prfrNgpolF
3lkLyeiB0DQultZCW5HsRnvmMBnwbEd3RQenAp1/wVGGoCQw5aINcaey7vVXY3ZY
kUXhBMVrbVuJ/n9npC1n7yK8XGu1wB7hmChKWE0vkNyWquCGfxo+36xsICYP3LEZ
TzQXXWHXyC+kjiDstT8ASGv2PxRdj1E+D4JBZwT4BJl3bKRl8tUxQMxtRuWfySDu
Oa3oA3LUR8pkSd5iY0Tuf+N3EmvEgIRsMFi5DcIjgkisLS/AMme4ciid2FzJOQse
xXgqy/fgylzibAZdiNo4vq7bgWsl3ORh5HYnx1LnK7rkJvRLkohRpCWpg6a6UyOg
I8iX+JEeDSW+kAdhmzCDgVFRHIJiySINeGCQG+JXm0a2u+Ey3PZ4rG5QJbaLpET7
l9UBd4eMZFcYavwiWwLgrgrpMR6Ql1VDRKO+XnDPzq+duB5YNgLdfaUVMSqx87NH
o2loJf/MX0y1dchWx0suf9UfG0L4yRCdZzyJJyomRWdZuO9LxNF0o3RoZbTGe6TW
yH6o2pyVY/7CIJ5n0PY5WTlEN4PGr+tWecVA03qPbWW1tf2G+loffpx5HE+dv0SB
NLA1iwMOm57bp7FwQjTLOmpQhsdBwWSQthLEvvK4Yqu14Se4lcejYKq2/YjPzq2d
AHSg0OSjMFLax8+E6DJoH3dwE8LniH0tlWNJO4jPxRjp4qIRhYgR/iOQGH7u8UQP
WMf9/CMELol1L6cktnRnJQ2OBYS/AKbdz7Ju/lvI7MkEhI7VxUE+uL/TxZCuDn/0
dIdt9Rk6DLSV15uKWT2E16aShAG4KtpgWKkOYBSoz683FwpULygWk4JWr25iZcBU
uvIC/52xLUXGBqCtVtLTupKsO5v80eFUk5ovgLe/SpB/e2f2y8sy7u8vC1eNiZ4E
gWeMoCBTcrzLNmtfV4qfOozrmb2PI0hJVh5D0g8Cta1IMl22A0bhac1fEHvs5mvn
w/ep4aa3ApsS7mzaOYpiy5pMNxA3ku43peGuYt6o5EWYWuwWfBZrQ3jl6RqW8OCw
yso2vwZEi7lMt1c+vxi2JJnDsH0rxH+o80NqJtIv73F+9tFM4AAEF3NVRq2jxroF
jrYicOzVnTmWinY+x6RSWj+19Ecyw++Zm/jZL6n9WfTcrSmMb0cAKsD0j/ebBeW5
5OXVs5Z3RHaC4p8u/3UwkmEEj0ncfpxFACM1L8EDmCqiq2Mv+pZv1iN/rFyctAz/
LWm9qU12WzkCI/zwb2FOpI4SNj1IRFj64sD7C3VRsZVv2tmBaRIFWzb0VzFKErsn
VDvbE21w1Ciyvou+RkKJzM0ePta6Ce2YzuCoSYpgJC42uXK/CioICEn7nIac8+Q6
9Z5pa2yjpvIdhtUDT+/z0z+lvlhkg74Vy6HdP3k7ZU2uDmQ5L3nx/BP6whOcKhz/
srZQQmvOxCpItyvWWE0rCzdWqCj8j03+ulMKwWTLpELPjapsPBRjJWJeANgzJfDi
6Tieh65UCjW9ddUmQYFtU5Epg7U9ZxMG2jwEiwy3G8hG7bN5kkKKxjB5fd8kbUaN
jxNgoqKkQxBZ+njCzFo2ASvHfnJyJTGsQK2Pw0G44NIzGZymPU7dQfzAiZlRjAke
cik3HdeAqC+uw51GrY63CfWKFtdlSVaqAOqQAxxjv03zXUjIVHm+OoQg+ENzkKz1
ttGEgjp2EDFEpZIvJXllhBmQ0H4ElGE/pcIy6dS5q17Ps3FVc72osa02OKztZZkD
o0ws62R2p5AJiJvKuJf/otTNzMBKsUqCQ+MhUs2IiN4nkmgEIC1gHsqZxm6XsPzx
t1dzBsoDuMn6H9oXUwuXftafLUwiFKTY4wJ2v5L4aeImWtQqll6tplPHtQ0+mCK5
8UfGfW/n7y5w0OhTCh+A1TI5SLEG0STynV/ue9O5Y3nl+jThbVysVR54u/4IMWuN
eDjDkoKDY90pbiyNfKmQuBl/5VxtpwoIv4FFBYI8OUQhvAUt6TGWAuB7qZtcRToJ
fykG7+VqYd27X2lfpRP+KTdVf9k5cwfCJNUuzL7ZhsvSQ7uGF8VyWqY6ZB94j8iZ
/HphKVSDwyEFmxGzhUNR0H3xrD21zbUMGrYYN9vY7wTM4JrA0U471JylB+UYWTiQ
Z0JunOa4UYKhh3KkbBmJ5nSmJizNF5h7pPrnHgWPRjp2CHavJYuwia1RAuv4isv3
VSE6tekJHQA0vGwtot95WrWWABDAGXlX/spKq/8oyL4+7ILlde0cHumS36FIFS4c
GSDfAl+G1ifdTkHnne6IWZflWy9AVj1/zSgagdrCHq94zfsuGzaytAN2Eh1vPjsQ
gnk9ErwJD853SgSHHj4b6+kCahXNRbBcI0tMhGnYcXN30joHa+6ztaxrSkRvUekd
wLEwaO1RDubcLqK7MA0qf69c8rxiibGgENYoFowb0MUfDLPh1R81AvZB9LE48rd0
WDLwe27ugjEy1VQgr8reHKJZAK1kYzivNa6DbQ3eFUW1lLE+NB7j+YQIsK3ixlVJ
ElIEOWwXwf6uDKutG7b+90cX5Bhf2rxXe8Meht/SYTqcH9Fbkx46N1hEXE6pXiX/
91uPvTujXNYb7mD+JxlZ/5HRj9xslER45wop01M/qg+dH7tkJIcKLYteJ1DiYJif
UzSSvzbJdVSAP+RceBnjIq9evCL6RYv+sGvZ8emiQlkVgcYv6un31OW9j2ERXeJe
IbNCt6SgRrUyNcM/ycJ4UgUXkJiFim6pMLJNodsXWlAxUpEAY1ZC+RpbdrtcHqGk
/I0/4Pcj1pEDHMexKOzTuH4+HJ+C4pXestF30S71AkkIFHDnip7wgYhdjvdBc1j9
8N0DC/IK+0l1SkwQaBdyuYHA5mFWGFIzWHR4aSkjnbW0Ye8rCLa++AhGpI4W+7qs
vFk6RAQCxy9yAJIz63t8/rY4snSuIEHNQh+3aeLobyPj3EOJoManJDDlwutokE9W
lAi7UeASp5YjbeFgHoztWsywnx5XIZLxSRibHGcRJj2PfCk/kDAEpGDyfc4b1MO4
+DWQJTf3D2lZPBVEVO6p4+udnKANpa1dMXCaH2/hqoukVJUsjW2Kc7bL2jtPm64L
vAFyPCGmGcecjIv9Yb/PNVC/FUj3dgMAGtiphqdEAeuooI8eb6OBQHxZJpgqQu/N
Wjp9LqBQV4RWE/VESNtbefFhCCepQq4g5HOjgluJJjRCmCNxFP/oK5PIfLfSLRY1
4t6/xJJnpDx/7P4AzO+ylwtDw4A/4YdvNVrcXC8eD+g26QSq/lV0DIdzWkfEyCgv
l099iMMUjgc3H1f5oflE+z+wE1D6IKlJ3T8j0KFEhcTcvG9VqZfdxUWnmGAHUNfB
Oq/yq8CQokt4eOR5ck1C3fs5duK6/uY8NRW8UicumJ4j1YeFloTyRpIzArnYfqmP
ycYpwCt/l09X9w+3qkVmIgyIkWHeRZ1I4dbhyfP9vvGmRDyEPd64besXVNgmOm5X
wuIUm3Sn7Kxlb5hFe05K6M3qbC14qeIpvKhq68iQCIDCSXxSq2gEkt+TqkCqxUdS
I7yhr6jp4TLZl2P+mdOqvRFhByH7AbBKOZhHaRZaI9fV9wgU5kngf3FHpAsCjHfs
1tZMzHqcncPpV/2HQvQA4AzMEOoAX2sUI2WQ5FzFoZzPxrLtpHZk1w0+uiU6n90O
/gtAqRVMd9aQ7aza0v1CjNLk2E2vzMtkSfyYFbxpk3nnd62uaofXSYknxg41dthH
Gzpt1QSTi3hNTuY5lZMJIknVh+sAp9ksVOFqlVjQ8zfHaWWf+xBwsFpkcCuLSRo3
kcSV43bT10IwsVDfSdu3yu82oXUu7avh1DaY88RtcxMMJ9eXrDa/JnT1UTIYioHB
nHXgRXDWCg9h7H5gmx7hB6YAvWRKPGQncHTdTiSirqrWF/TlmW0le0Wg7tBgPi1G
i3sms6F91RwBdGwUF454LEFl5bkj4Fug/Chb4uaEsyZXQFYdk0eLU2rH/vwfyW2l
XF4J6NOqYycSSFKxV9hc3xuTaoLqr5wPUPMV+hV5nEBSUt7KSUyfH1i5eEBiBKK6
iReJf4J+cmf/zWor4isCC14fSa5qGBHN5HVtaUsYaMzpj/BJH68Yv/MTI3kcIHXW
uEQ4Ft5IZEWhyK9zoaxKMj6F5sMhkJlvCJXJL65AFK2u0eQ3C8hZUYG7pqD6t2a1
l3cNI0vncmA/RuxxPFf7YUf/R3ffTYlJMraXzcDUPALVYSpafk5KhuGpb5HuMbQI
61ETl2H3JHQvdLG1TA22X7qHdMuIwVi0yu6vGfpQbnSiqrTcC4DC0VYwpPTkktP6
EFVoweihLXMfPUBtJ6IUmb1paYcKQXm6chRSS6mw7gxGB9CqcMnftnObR5ATPLmw
SteC96VfjJdfcOwREOCCkdmkZXhi1QvNs8Qx1FWPwru27gTblFq6HLIZqMuxpKyy
rPqjl5YIRjBRkkkyFToqJ/hnxvOQKdLluj7IxsHujEL/sO0KCyHFv3va6rKyDl7t
mYlyJCVpQ4M9TpmmSnJFe39nqxyjyYGHxLwBAYZ0jfGC1tPCwAt6+VvgP1eYyR8/
xMPcrJ4tisQXmzKGqp3rpYNCutt88CxfhCOXF71MH5nOV+qvS25iniTfGdDoKrMB
oKDh4d9B45WWsgfjKiGeEBBo30LFahZ/jDaZ9rNEcywaWDp+1ZuAfP5hyN4+uFOL
Nw/2nF7vnw9+PzzRyqmMcIHRcQBX+WPdOaFST3IOFCCnu06rgend5qZTvOIgHcaA
nGFacQiwWyv6C6m1nuTmbWvxF+whsXjTxYY6w7PpRF4o0xQmu9Gz1rvKASXGFTXL
+Vefa5sS2/pMpH89FqBcK+WzMICK8inglCZqFmladsMSxpesG+PrtE1DUEr+A7DN
3Uuwa/545u/UIpBcuFwAhqJ/nSmrNqFDdTPS6S/TuuMjTnk8cUFtFwHpSM0nlqbD
wyYX7nTLqeHNJBSELg5RDPV/Uk6akbyYfxB1OUVd2Mc8R2cqEKmk9FoP+dE8G3oI
3s6gEPKp8jxr1r1K61hAQdXDlAJuwj1lJAs+BnuSnO7i6jGZr3eiVNtDWFlfhLFw
yyj/I92VkQFQmgXaHzxrsHw10b5L5KX2XsWmrDtzLIK3MmsNN10mSwAI+HA15GiJ
BcCu1Qv7dqZNGnbNSdsj514F7H6eDOkHuPOtbA4vVnx3xOR7WLYD22hqzWriqLEU
VoU3SlFzWYLS+B3FVHQWqnXM4A+oORyiuFTzJ3JauXdZJCE6Q56Mk4bnBBhSeBWE
Q8Pf6qhEz3WW1MqumGwzCpLMnBcXwHiKEbtVLxqYB+nFuO9Gd33+3awbVIUOoIk/
m5qESvZFILQ9xSZ46lmYUhoIAnvcURe9nzigVWt/tKHAaeTKbmwmrTfpGrCgcJJi
Vy+rL0pXuEboet2Y001Q2OPwXNXH3R+BVjQ182lqaMTiKor2mCp/B2jLdCU3Z+Op
z9RAESsvgYzR0ydKrSwm83ET6N38cQQV3a2uiD/ZRYX6NbWrpsmMqksIqdjfXZCN
XYNoBRlG5cBp/mCW62oOwTx/XEzhYWEj73ns/w5afFzDRAeW+IsWitvSSUtIw3Im
XOnxk8AKrX+4+ljPMlJfcHBMeB7VVcIns/newUtjiHb7mkjgloL778KzPPwY5PE4
ZudPk2ATTYHbqouwyFu9a5uKIw+yHO5S5F37SY8UlxaQBok888QoUbfKOTpW7IP+
GlyxLJID8YWY7YLWCBNg0qZG7KI4ydiQFP+ySS9f3nkj5E+q7vtKWYlKa5m6iAIr
nKHKynDt4/lue8pQiAu4ILZlPSjPkBYn7P/KPjVyM50sPTo49MwvcWUDtDRWD+m/
QRMgPFliaV+AIhk3zDhJPKoVuKQEa+JL2plPk2lBhZxtBifoiKQd/hYNTO4a0E6f
V3SAoM0KpCqQ6gy2X2rop5W0PV/hzzaPHX+wPtidoQDhO3C5h2e7CmYLsFS0EYhS
ztxeY/3+NrnWcWN4iygrsMtTruvI2movY83ffEXQgqzcrY/VvGoBzNYyRLcg4N7+
ei3ddJRz+4AM7hIltrzkz+nsnk0UOzm2tt7ZDB1UukdNsL35M7F7zuto56BDZEAE
OX5DRy+HYGg0YEi2BAFuHj2HndEsT7ZCor50ZeQoARpVXzfXBqmDAnv1vCnmODl/
NMGlMadJk14v6wqkhM0UlGxUD2X4UJpq81swZTIwuncxpoB+tx2kWqKn7UaQCoHN
ENqUyan0Smdf61bNzcORMY/j2VlEjWz6cL8FIEqV7ve6YFeJQshU0voP/trOe3yu
lcTG1LiROzDcdRD38SofuKqGJhBqG83JhgSDHWG3jMYB+uJVcvFPLZZpRaGJ/Nei
/wLqiRVYv50SP30II2vt7lMVMwcvNJB8nHTbbW9PSQuK/k0S7NAmC6DiKunj3+i5
YEXe/b7cFGxk20q8WdzxlsdkRHCPW2FBRwHV7Gg1ntVt84BeHrIVBM4zuoJ7tTVB
9EL3D6phwk7EFfEu7Fil5MCNGR2wqEndZlUt0hnh/9haboifM5PqHAgIyAh53MKi
i3WL7GAOBToT80j816aUkb+5vZWGTax1OwKkXJin7OJdrAbp5nobzLngFkftrWU/
5DPdBoGjJMRZa8QwLTNt82EnqvqiTPB7mcAELUFLFTnmMcr+fZGkYCaOD0oCmzdr
cQNmIi02+cicuTaszcuEbgW1wcjoenJ8GNsXUXTxLPZ71fP4wOKQ73wyHZBt03Az
LlynhUUsIT0uFVz3cqQpnNb63egEr7ZTwfFHTkMrSzOrXWQF9iOTJJ478uCF2BOO
h9eDmgHlN9n+x+8sQJ/5NWbEE4t9r/Dr5IJC0tVlpxMdS2qwlp/1T39IEw81tpau
TAPyei7ZmLdFo/Tpvt5qEncL3GDuMjRU8SQrf18Upnxa6SAS9AUGn1nK+dGh9Mxn
FTXEYnHMfV0Qh8tClAbkckpNyTyApvg8ozOSrfq6UIzJ2CkzN3ul38NOzJHSQlFX
wYZlXuR5WSQPp5L/tGJ4GI6Cx7U4ouFT43C1uYUhgnYgdTxWobu55D9if7/3SCjc
3WGiBjB9naUj/HUUqa13UadDR13uQNeIY0ppVkq2lyIvnIv+OZwQl6qjDT75F31r
SBikX2rp1qahluI6aGIcyXCWmdPgUhxcMOTYTRYolOqewIxzQwkFmh6f6FVj17F9
dsWYgOV4oFddPS9ly2vS5/ii6zZcVv2QVAokwXtvGd+ddO+JpeapbIcfzjLLQvGI
FRmDocJq1NwD1dXyq5AIR4TbAJ55yZtH/kU3Aan6kj+66AUqdF8IR4c5nEy8LqP3
cuqyGJMjoW8kpaQ6DY5a2YWPXcZ4MPdCRR0PKikCYromMv1q8em8ITu3u3OYVnnG
wwx8/sKcJvKzyWShAX7ZpJCVI4qI0JtGA8JdXbQp2An40vcoVFYIWqCY1GKCmLQ4
jvoHnpgPrKnmqecVWIUPaSXgCxoK5Ul+GiWoOZfHc0qRtqduDNvuhCryMccOcekZ
3cnH5zwrvE9nTrpcTzjQJFGSpOoFDG3CN9qD2VsvECk1AHr/uYas95nlKBghpgaX
3Gy4jpl0eRxlpjRb4VZ3pWrnMrjKwhDMn8YZnjQJ4JNScLBX7VUN5V7bNv+ZKhPC
9y7UIb+UPwNzw1lU/ox5i1FeqMAXsUJczN0b3qKYQpxQWZSgLqriUJtDWSCd/kk3
/pbX6Z+yYBF7jSu+m4KycK22iWfD5Y11vOMsLNC136fiMnubTkK2lmcnsuVw1Dr6
xuzLMORCWngjPZmQqr8VWBKI3RYWjZAWIpHSrXPZiB/b7CtoHwPcVBGmew6ettLZ
kbpWMlchzFzAMzY+8ENtTuWvcqrJ8jrn5EReFJWsAtqw79UqxyyDV6iUN9duiPW0
FUzKt0bhlafC+JphQtz62pjlctdCYH5Q9UQ9ynIf8nbkHG/TNbml/IRTInO0yUVU
lyELzf9SQ/CfwKRnqhgBL1segugz26u/bTTPQrM9C4+JvNqU5POlMei/NIEOT8iJ
gwn6qbwUScsTE8kcMYd7SJW77Ypcd05+Pelk77DnJ3xMD9aDlMyHDc5KaijX+e7s
IgbF4XIGrQXMVUtPuTJy/+lfK0TEh4rArEA8H7SgSvsmu3X8y42E1I5M7CCXd7ll
wF6cWc6sWGbPGmd4VN7DKLKXJeZdT6XHGCFE5czH3un+zSqk5nMjtvC5ha3SJkJN
faz83j9EFShv/1n026qmLNhC96SM/lZst7jI58lCVRzieBxaxEX93fOU/Aolm+I6
fKvowDQHwHmCJs4Ub6ux16/HJSuuzPjEkJWEK4dV+J8RR0tG8zihs2WbdGOcQvmO
C1pHCfAOwRlfe2BnkZ/lR7bgg2IEF7dD/esRaMTwebpFTHGwsBrpg06gjaUPuUp6
HOwtQGFxTKDcbSzLI8Hg2jmBTNWSiixBiLJtMuSBMvM4790nMoasuMJF9OX604oX
FIrmNvtXsO9G/f/ZtL6bvxg7n5gzadfOYsTxPVSqNHq5IL9dzeTuESOBxMi3b3QW
FEOe4TdiHbNe8vQ1iPu7a5L0TRL5fTLIARgjz+t39oHzjAiJVGLZ9ve3Y+NBOcaT
7CG14w7ZfAvJpmqcO5fM/S76hvfbEeV13Au2UBfft12ZE3sWi0aYAWs4+lRQCCju
+LFyiFXCShsy/clkEqeJkVQRO+0uhsTnbLN/ZsDqVj8KyMnvRBbIlDUUPnCo+oHP
JUcRketVcH3K12GNrBvu1dp49yOJV0V5pB4RhmOASN/eAbXw7dIbFhJld5qXowfT
L/lLoAL8r+YVNDTiLQjIm8yGlZDvHfCtzFp3GsFbb4Fd36NuW2hDhcVjCg2utG3T
3NAB2JNBtmnaxB4t6j0JQf8YtCC8hTZBp3nj4I19bfgZfL+zx4N5mxzEuhFwReMU
I9EBJneTh41P1I/MMMy+C+1EABaJEWsJ9HG9gjk99dVcBBXkiXMWYDDtGkPgf9Fc
gfFUKKVLVHwUGUC+1AsmzJ+ZcJ9OpJfbjkNj/jf3j04Pj06Il4XXkPE0+c/OI/B4
j8rX/v6JMvE3HvjH3vmSuTqe0kK5YKmz1xgG1/L5iMzURJVV4d2igKw3AEvxnvEV
zduqQqSKYLUNYbAOkNXiFIv7Q8ez/Z8/M2z0eLB2xOPBeBXd2XKOqojP5uM7P2JN
InsiNNHCMdimObhW+HM9xwBh9b6HqBV227YOVtW4ruaNS/aDWJIwq2WLFNxirqpf
2G3ftczOvUudpcOGKb/kN0cIun8D/Bj0FhvBS/zJdhr3lHKnzZj1REcBWu9b0TGb
nohS5fxOgq1aU7tXsh0HpFadBopJoseHbu1JCor/UoRnGyQWdGE6bs1oCCqDk2Ee
+PsNE/7mtXCAxPLaKDrI8zOWrIQXMa/gXV+E1EKNwC8QaM7YsNZYLC3Ausqzs5mZ
Bhqh1sAHEnaIQ427NmFf9BU/gajViGVi3Jj3+Q5fMvh75DAiLH9N3Kg3nscqc/z6
3wfqkdYRL/M8I6bqct43ldgjW1/Hd7Fa1M/jb9f40W/9G3igyMkqv/Ed46FwVBVr
49HrtLfAMQgdYpB7dJst5R9RAWyaX8YbEGc8HfBO3LQNTzACUzzk9IV7VE69RHzF
6/qs1Mi57sVq98wjoObWRFbsoi5auMEazzx77yXVcuoqRJRlRsv5sqekpOATFCKw
wcYW+xxbjEKf3Om48+KeZ9ssuJiFt4v+SiwhwVvMtozyg1m2A30stbq9hRZFQLxs
PC1uHMu+ykeYhxPgpz8A122QkSfGRSBp3tsnNWvwS0cmU4HU2n3Of1+YNqlPqD8y
urNM4O/xl8H6nPKNYjjY2YJt5CjFQEj2W/2XvLMkU5Pey/tx+yaHRQCzslAENFJ/
Sp0Ks4u3H99Kk12yTy+WUl382c9d2mQYMImRUD7JbDHF+PqninTlk8U1Twf4DJ+R
P+GlMHDAhhIebNXzt+J1F7mKriLbxEMXasHySHsNUcxPhh0E3ttvnbFxiPm4NoAG
FHboBWJHQpwE6V36J7foiKASMXLtZlqS9bg6dmVh3FqQPkUjcZx2IbaONK5MP5Gx
2ZJ99ydN+qcSbMqFFy0cha78FQURS9JLcwBSCGxrkCyX4T5ro6SVkNCR3Pm0YQYK
4mLtOgMHGGWFbhsC8FeTiBxdu/Z1mTuFHt2URv2unS6vvHXGsQFwDoydSULHdRJ9
G+a9RsnDHx4PbxW6asZCRppbg+x0kyb/NoKFql/EN1wBmYoUL7tvMLlUXe3Bwx8o
DPZdTKRB/zr68Ug7zhOx8iy4Mq6EUa2/XvWPcPoU0tOKwegeX4wRfPEkjuHW5XVq
Nkuo6aUzP0U6L6I2jL55fMnQn2euCybzGhsEJq5MXzPt1OzlCYt9wlqztIRHRbFD
+xC1t4JFzDmWN9l3+SSbJItv9GbwXDz119HJBjpLrdQoxp0/hMfAGkP3RcoyhztI
iCa2zK6Jda7jNG5mU6HLAEa8XYZlUbUkmjjcT/N62eLM61g4/n9OWczCHfKRfE0X
VWbBn7V5QRlPP2NR5kBkkvZTYxxbl8eq/Toi8wUFeqgo6KYf2o8/kDGXm1R37UxH
KXmSzNw0rNEu+XkBI7PHR4B28qhimICDbRjMEPQHVQiXzv+zcfBrK6X6xmzSEiSQ
ggGTIeWPRie1Rh1CxyyLxcp2C4AdRd4nlYvKrPB27go/o7HtApJAWZLTjAXtTFa3
kwgdjbwsSRRUUesJAaY0XxyAL+3xHgZOxtWQKoT5SIuNoAsCu4a/VUla9ue/c/Br
EFEU4xGsmVxlg+E4Cfutj3zr459yxcb48/f1eIPZjSB5sJeQ5uJ/66whSO77eYSL
sP/0ifIrPEZAi4mdxsKSQlYmAD4t8Wy8BRyZ9F7B90AWi3kCuVad+L1FQ0cU/f5p
lvbyx3szz0P/EVMaqmQxh49ERDugJX174fn5Q4lBX7nm8A7OZtaIN6BwaphlxHE8
d9204EI0GLUNKhy7ATtpMRXreISRzSTYKsoOmSUzxGC6Dl8CCG/xmbInGwmx1xKN
9gkIV3C1ccqhHhdb3bKc5W07fzJykAemHRADr2mu83Pf4oywwccTGIbjhfbPST9e
G1nMdDRclczCwN+lh0pSQhPz+Nzy5q+HELJpS9rKIXqISSq7qAKnd2zz8TVoskKx
TSGTGeu1wVId6GxgFqYCDhJYa0UMzt7EhB97nAzkpaJMWv+TwAFeVJAke2XXe1HZ
m1N3OjC+ZgToHqjoMMwhC0qL4Mp4L5AXOnaxgA0V0rLiyUPucn4/B4ufvZ4voK7S
mvfPAwrufBgcAM06ETM1L3dlV7jCh26GljWYLgbgOHpFbjBgoDD6LLWwGXKbjZJp
hBGxcRQFyVB4BKinNRvgcK1mMPb3XkIII6M9t4Ld+zcHaWVBFk1cF7FhfwrSFYtL
u8yhUCnIAllT131DTrmPwsmHFMsHJq8vjNzn1ErdVBN2wNVjeriHhXjAtrkcpeL9
BhQmViXBEMZk3WJjk+7OLvKjt9vCB2CJnnChS/2IxuSwBczH6iCXt+QsoKSJfuNT
OMziRZqszXVzk4SEHE6W/famdgkZoCt+oBd/9gVFLOO09ZC6n4S1zNFGre0sg1/N
GWqATV+u1YoJfI6eaC1Gk+P/NZg8s0TSLOS8hyV/02SrCFrUmyHUqFi6dZWdcoz5
ZNplzDsuHHJvNVKIsKDOmqcrVDfVsnj+VIWFQJygAVauO4NdZ4nEvXDuAAZHc3Il
Hn3SWvykTemNkddnxUvB9Jzp9fEH2pM7R2G5Cs+sT1uNd5lG5Oe9tmUt55jTDgKZ
VdSSTcFIIGuEdUFBcqhsI5I13Y/cY6JSiUPPzom2g8y77etgtIjWJ4hLdQnEpKFD
CYV8sZ5wV0rBmB2/gI0XGXNtivUf4NJxiR3EpofJuPF5Qt6Lz1rg6gUkWiDDyNeV
zbGK+TRPy/S8/vbWgQmk2wkWxIqvwOMh4lqDq/zMTfkQMbKg2+M/c+y2wWb8mkr4
DjMRgE0JhMIIPejKua8XLdR9Xz+zKiBIkNtQSYkmluuJqfADExuPQzgR4qJ76LTv
hd+jNWxwCxQ+ac3dqoSjwdBX+Ekoa0uhfeinMUa3CVRy2tTNJDiJUMDSyumLvEUs
elx/o9RD4i4Vg4tmhlr2G+CC8lOz8FkSYbkSV4x3Bc89Mv2XnSBohkwgI4vGv1kT
+Jsl2fZLeycvKOyyr7T79pDxhvh9GoAFuVtUKVmj29srRlMXclv2hMDrfiqY9Zp3
b7697c/I4ADsjV4DR5H6ry/YCE1pEesAWY06GtQ+ypeE7wdaYwY6pWZyelfuBBZr
SUUzjyTwS0W3YrCyfFEr/i033zmzqOC8AMkniCemNXfrgn/aeUkZlfkh9LJwdEsE
HnAz7QxQk9rse10+4dWsoTnFsWDq8WLkStQ2ugEvzLvbvRXZ7pfk2Aa86fgWqVse
qOB8gxedYCc/bIGMTWNdAcWxisBvQCaqpnFA9X+6H+dcO98WLk+BFkiUP4At10L4
HprGbQyCdwIzdKTZJSqYjvP7hQeuU4U1ksKjYwE2/5LRmcPW2Ln6R1Q+bf6MtG33
kiFKzcaSVpmGG3EtD5BcyuBmELD+Hh/ZkebuIwkMSkPfo1f+RebeAdCeesRKBu0d
UDdnnNguc2xBDTBdwMkGV1qGn7wUmwOEqnZvpxPPygBmePflGzKqdDVqgvn49prr
qJMOuq0ciSBEZpoMc8JFxJZPC5Nd+IE6m7sGBMLpBWkpi1Jw45FycF8jsplMI/Tr
8hwJALXCjaG53iGwl4TbiBj3Swq7joC7v3nzsYENUimGb51ldiAu1GaRkBXLcG4/
wqCE+nBeNIdgnEeKRZ9RwBSHyTUx2go5WOTLFV7oB2bYldqA8HWXTasfdlmS2+0d
YyGFZZaow7hNAA9HCw88SVxMrqCmSXx4363JNNhC0bk9IPBtAFnHY/ODBOZpXeMx
9Fa9w1d+Hy2c5cxceaTXx1OLmWvp28E22BWazldfcd5urEghQcOjj9PetUlo85pY
gkxcLkUGX3FgB5/QK4bBm9F9XZZo07icuPxMT3LLLezFU6a63cQPsfMRF03xaq7x
HuordW2RJNy0DlKsS/pNYQbocFQvShdbpRIZ/QM2vpGUnp6/gkbRjDfkX57JUhzE
r/iWgh/JhHPFPIo73LTHwJlW0+JSxWyEVSZKg4hJdCv9v42KZNatlfDJ+5c8p9xg
Tj7J7Z/wjvV8h7MikhqIjD9i5f9Xch7lAg/CsakmxiROvhgdBZ+Ju/HsT3ohGOTD
ZaVN5Q0PNXDc8K8X0LF8bAxOP+8DTIfUEVNFxmbOxubGKkXtvDwR6kqqqk2d0BUD
uyvUIQFiF5twAI431twQpjEWvW3pBEgFf+biIb44kYvb3MmJGHVagT6YGb8GJn7m
k5xLsW8qQJlr41AhdGHgqYsL+UvBZznwqMTFMFzR4SRzylYnyPmx79Qa0vR+r8e+
ORCINPC3QpIHCYtB+T1UVT3JlXRQ+XjJzAcme1lx31npYurcxtwgZxdY7xnGAvdq
qLPT4dWyyLhAXj6I6QlToVthurM7bzpYCYy+HFvpWSBgnW/QJvdWq35rJi9HOlyb
sDcYRBW9cxMX1NS7ScoaJ/CsQYwwtMFS0t5/5yHGqtdXmfJb00/Mg0PaldSJW1M9
w+J9jf9P0kfyfy5XOsW/3CmMFQIIOCpM5DHn86+fWjo4xqrS9giWtVrad7p74B3d
OC1DbuE1EdL2HwEbXo+kHQ2lLnRwzJxNMQ03VmHtr87v1/hWLhnsLcFRo5JVLfWz
ls0YxJy4DomHXikpxBuVkSRPf/nJ0mjbgY0YX2xgUhLNFRNvLYnGf4vX7lxZK3md
MzgufMEV0NuFWup16yb0zPuC53s5H3hW3fmUsnQGvo96Z7uToa6obcDCz55r1vnf
VYPo1QSjgFUZ4MyCRTNS6ZMymIBd588IPW0vL8ov1e1/UyY9fjTPbYHKBjxNZohj
JZauw+Y9FvOwdyZacjtQgZAzPaIrELwCeRxfrojmBpe1VHzKnBrMGcL4X7OfrAi5
2ejyD/PTbmKdgJJ2uakHhHIVloGbH4bN8ydVk0K9hE3xmoh75eZPWz9v2SvpVndV
iGQuwMgAX4hHcz/Gd/058PnJuxRMpsa0Sr9rVHZGnmmkIhWgrCWPqBOcDoCvH7Lb
+weEBXRzo0olxRt+dhS20zKffyTB5Ff5Ax7yOqB/FMc3e+CdPFU1BFVdccWMP1H0
llFgsYgOq1S7QtRTEy5g5MUOrAT2ld6deHrK6nuXZj+KLNE20c1gJkREyoOvT4NI
ILQqLxWlO8cMpdtXCNsKZ0pVqca4Ht8fYPw0UXuLwlhmEnkv4AER2+g8YBnr8HG9
3TRaFa/Z7pOAWxAKDyLXSn+/jK1vTznQpP3qrQTRFj6gvza02QozsZNVU0rNHOjd
uA2jLhnMZKTiiar6AOkxhG+j3GQO1cX8PZVv2TW0CayB+Lo/ikx0SqVoFIxWngLu
Kdd4BF4Z+lcHw/kNgPU4JgG5cnzeLTJgPE5nRadoxk4s/JtYowK8ikXGVvnkqWD7
4aq71GkrapJfL+Tj4Yy/aN50ZddXGQ88w9rj/IZYjHTREyKNH3Gj9AgLYBA+kMS5
fHfR8o98fQ5EpKIjtMFlQdEcPKpGPzb1aHAUgccg/0AF6t4XIIXrjfCjGn2iU+ZR
/Nrb3sxVfNcrHDrx5PR41Jv9N+yk8xIzrRq4m2XzVMGrZhJZb0yj4YwyhCUjpSHV
ScvUSpcUSklKutAnAcTNNBR8Essddb2jzUPPyYZRps8=
`pragma protect end_protected
