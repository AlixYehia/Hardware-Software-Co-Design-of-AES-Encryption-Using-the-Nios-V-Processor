`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sL1khb1nCrYUU7NUXcVZV9woWobrCAgZnLagOVJDcu14ArAaBQFg3a6i6d7PVDI8
ax4kRlvYRx8c7cKXKWhTAf8LSd5VucSYyYy47R1YeihpwA0ylXqEw97Gy1/YDJ6d
4QHREQBZAzejHBK/TYIIrEH4LwSftyaiHKbXsooE/Ug=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10032)
2Lv7Ichc8K/4n78lhhNM8VypR7jAGSiIgM/XicCboM+IocnHz4qupAyUYffO8MDu
AecJ7HWY419jHXz7iZ8v9jSQA81z/bVBxHUH3xI80XLXOcJYlaA5/7FefN8PGfsv
JVn5FHM9ewXskgYnbULnxFz863ZcHalijEDAwtu1lEI8N2cCX+Z2tLLtcEWcZxWq
lrrZl3u5oAZolb1gMf1/IGFOq2m5/R4nQb3uOc+UPYu1ra+w4pNIq33WCisQF68P
lW5yQwGopaLQascJoylPxaKasj62CtOHLbbDHWLXvA47DJAL1FM9wTKO1HCjI5wa
bI1PGJJwifTmnnIRPqVYbdLUoqaiXiS2OpGfz6eoZRncVh5ooi7wxQqU9vVu8ryg
v8YyEaqGF1Vt7aNFI0OKojvjp25UR24EbEc8gmorH7iwSEQq0PRA6cA4yIBH4zz1
U7t+/H7sczjnYizyU0nY4ZwwYmi8MDC7H+hj59hrqyko+jUzmbH8LM2vhWvNgbov
9TLRzaR1HxDv9LndP2wQx9vMh7mXzMZQPj8oqCr4F8ImpML6gmKbXNGzuvhriroB
ohdCv6k1Dm+9BbVw20lhlUkUFNam/KiTYhgdLMCDZ/ohk7sLcK6F+nR3UJoykWb+
diPsuYRM+qat1sFxPQfBgydMdZmYVL/Vt+RO2uI9a2gJkJL6cXSeJU29fPjyCxsy
gdyEIlVlC3l+d7wUfj5FvxBdrPbOFMhUw47MIX9EOELbAFIgzzN1SbIc72VneZTc
Pmrun4DHPCsyJkyj9ST8Qdkw15SH65BZ2sBIAe0oUQAkB/XZrNgz2hT0KK7ihORp
4PHGDSJHX1fLvPBDFs2Rbn/Wu/62H56CGI+XyFYEIWcoUM/sPsMpFllq/A1UlDRc
hoMpoBuPVwSKU62K9YTStQLDWKpO8kw2u+uKZNdN58uOTv96WsXv5w1UhnDswdEO
ohBhzU+JovnwHVIXX6sWJ67qua6FhXsVlnqMCB4gRkUIzlLpYTThUmqKvlXsURHh
lwNeE9tcZH7E7QENHKkx8KHKs5Zbvy8+PcNXcNCxFH8hbq9eH+jaqTvTak4N6QMP
W/XxFCfA2dIGJ3zzWpdy78WvIEIAMOEe+m2TXMb+7oBijxVLCF2y1CvCBl8z/5oy
YxdayFBPgzaxQRxbNLa115RbqyQxhA1E7bPZ7QY9yFxPGrS76xffHCNiwJF/SeCx
lQAXzoGmHX2eNyjd2AZ9CAXc26X2WzvCFvocYvV31A+hYunxPsRZ/hPgvkMRJatU
j+v2J8Rtt7FHFRTpVUmfRATOonPmyIQ3gcE4tS3l9aE8NGN7K8hqK9B1AoFfkVeq
J4E/t3+Xy/PlFsp8fnb4TtPe8Z3YjuTYWq1uCeh9MacFoaPdgHEa7vWYfnURvOUw
w4ywmWr89GXrbIdJyKqDu/eczZTZUQEWTDJmpUDiXPzLzsNnAzzXCjjoaJvbAPbu
s2yKmJTj4ALPQnRmw7vUOWl5M8VsCFLr7hTwv6S9kDmO95xHbLRr+XtxeYLS9+yP
/YR+2jSULkIdgDJr/I7sW4Q6VLMGQmFiHd6uVdQpUyetOid/e6XHBlj7IQjgkfBj
NCJKjoArWhQzXnwcb06kyzXmvQII8VeQfcmnVY0kwEB+mGJ0Fs0+We0B+c3DCHr2
1capM1tqXbeIt4WLWslr8sISsMkYEIUPnxltFq2YcjmB6EXailuOhsKUu1eZvpNp
x3c0NmBY55WfX8XtLlG1rt7gHMoEBeKmJmgWKaERk4Wyy1Mbh1v9y/Mou/EKaJ0m
q4BT/YKluJ0yr1ec/iHeR8CgnJa9IDFfIS0UElfhI4BO6BuRt+KcsZS//9UfKQGk
TZd0eDpG+X6AGMHxm5lxJcY1AAvu0t9+q2tku3POWLo70+3Qx80DyrQjPylyXg+c
WumFSZkCgGAJHNSpOAB/GDCAZTGZLuu8+9vi9xdZ1f3CshM61Au3o5qkucW6vift
wcW8XXIX96F7jW7WhkUhjY3DOEJslBYbMTqmruIEGgfuhObl/R9YDGKiqgX1nZa5
I5C6P9bfAA5DZXTvmXMNMuJNeOVfA6q9wUzoosCtFJWHuboDejk870UCseJtAPaG
PDV9Eu8FwhbWheoprCRL76oy07och6peliNozEwVlitIfmAiogu/ppoNDqsyoaA3
BMz0Tp9nfCX/L6GSlKVGg89wlDCicnWDyXCR+/4CiDNX0c0uHy4X+QfAl9YeV7Qy
Z5WmTR0CDCiCbbvIPx2kz/jpz0g/s3bWPbvDA+IkN6TCkEs0MhFBPcURvkHWdKX5
WPCMq0SqzBDAOPFYqmFvAjzLXeG9v9X0iHMu9b1CieiPXC3G/2RUyBBtezzJw6yV
cS2rj9U60G52zAJJ/mOhgKYP1TashAaaz/Mo79++12xH6Kh9iBkeIxalXiKZlK78
ylbZIOGK0aohoQi8pHsQ1HnMeHpKA1FAW9d6ADug3uiS+bjTdYe/7g10OMbBmkdG
U3Y0/2L0YWuU9vQYXk72nokvcYwwH7LQ/vUcrzJugOr7ZYssBGvaAZp14V7TWeoN
CCI3mqXnVOQQHXpeSINKvz6s6g+waWDyuXZ+lrNLO1MSCeL950ezD4wQsjszn8r/
B5xXLjoOXnEbpFc4bY0AQGqX+ML2ZhBzScdd2z5QPTdWRxCQVLZFYSPdd13EQ0EQ
4H9/VRXECtrhSZlrRusVlRfN9jqWIFufT7pCg2oLVTGXyDYFtRubSBdh4VpsWM4i
Bp8nGANX4V4a4pfWVvGhduelVElXa5TJDfU59Mb+gLFQjAMuLHgLHuutMh+FPjBT
xcEBDvVY2BtiHAjFM73FNaGaPO5QjqyPuEQvBEJotVI0qmJnYMQPWFmxrSusmaAB
UrU8eN2TLMgz+9pOSQfoHVb9csq8p6uVW9WzBC9jjpYNOOKmPNzm42pYVAbdtDG8
AAZhZO3cOD4o15Bz4HR1EgU4HkqPjSrg40A/nBPDbfpLCaQHmdy7c8nJOqWooyhs
eLE6bZsBBvL9P1hJYTBMiyD0MIB00ohFHsD0GMwJ8bvzpgt+ISRhoms7nWtjDluu
aMDcYYTiZeIxHB5KpZXKYc9ZZ10y2vDf4gQ8fkQSbXnWKcGrxD+1VK1osSwkKNLX
UrfmZENtqjX27tyKrsocYI6cAf4okKEVwjBxHh3gojMRWyVz+21iaPSyOcV0jtr6
de8p5mzHwRqA01aAL8wCLKrTBRUv/BB/+fkjsGD6oQqJW0NwbKhVThd2ON4KWrsq
5dmx4gsy1XTcH4/eofEl5sCRMB68jEkU564ZE0AXwsLHWjfkvuH6WqtJJCRaaHFz
J628+EdvLSWnzOpbKbOOZC8nRFLD4BWD4HfD7hBhOR+fvSX8jrUx/AYg6GvvnyM4
ozi1WfCDNz/zVEfbU51wPAQIPjSCxAKq0EYKJHZSMKMa9WAy5dDKXMO78KLLHY0h
uhBIqoFNjAR+qtNUBAl8pUKZHevEL29c7jtZjdpYgqVoGWIMFNF8agH1Dc1u6/Vx
sTkbFSDyqvUgUYig1leMM3qcjBIlhKLw5N49PN7MSy90ai23e7GH71kx2t98HKmg
O3FhOEeFiBrBZgUJrmzmBBYqijOh2lu37kFqJDppZLj/W6SgA+d1hGoy4dLMD18J
nc/ZWjBcfN7LB9X1tn+Vzw0hvukJ+xLGIk8WpLa4qEUbWvMUJ7ru5kgBe6zVy6pO
RBDFwWJUMr9bMlyp3JIK++CB7r/nnCxDE+EQVX1zJO/mtaSQmcgt/rIcjXQO4EoX
A78n1vxBONmMypuYBQf+J5Ueh5VqOm6/R8NLgB18YOBc3cZDvqBOgwUKpRDCqGbm
zACVJGpm4LwGaIsfIsOouJEdRrbB/APSBsEaUqSgH9be4dG1OnbOVgZJ6d2Zgtoc
9ENdjhxbKQp1Aus7jEwjbov/S5KOziP3oryfBKcNwgsfpVkDuORDtO43wRkLdkR+
ESK6PJ35YoiZt0wq3mJVRHBtVxCkO1zwx2y+yZyVn3JSqYDoqvdz1PQ48KlMjGPa
nHxcVVLcEniLr9BcPSpZ1Q4FNqZIqEY5YgRIH6hM7w0mVXVQbcO5/yCcdxJFlbnM
feP8vbB1adeoLRlv/pH47RK5UUhbMvLHhwzqLkcqxICtdUI6FDdEm1FWAeAvfhtS
jUecFem+Phyxn/+PXtr10y6R98+YyS/p3qt6r7jglmZo3BG6xeJpDRQ+I1pUT8kI
4Pulcb110BCnsfXY1PAHsbVTW7NhDGE/GVz/dW0PcnWhexK0IJnLx7bOoI2Qmuzc
fBYHX5Y9cC2XJFPaFahbujkAeSea78iMQMudrW3XDGyQo5SiPSw67KulDKDuJDq+
YZIe9YiF5U2T/GdqMcRedRojhHovsfXgHAk1nF2K3KSqti+7PMbmyxYN34bMbyIG
6mbT1pqTqI1igXFjOwxMJzHMESa76Va57UuRJ4PsCtjilfsTuh0BGzexshSIT7y6
7dizsGoACPBZR+XWfEmRfTY40V7Rksqysr3cFpz5KaLP6kbbO0TL4qXmzv+M349H
WzC93JIcPgLo8nIC29CkEZE7PbCXq1dspsf6nLXER/KxCKzLQ6o0J0UVDm4IcM2B
BD1RswMDbjOm5TJTYquazNRBi69hTtE7FjQXD1Jxe3PzbLox1W/ZaqYX9lqKyo48
MRbFeZomOeQKzo3a/mmHWyv/ox6pHoXVAvw3m1JH0jr0+hEjNJCClc24bgZgrAfI
uqFTHYgFNovPz2/bnXIDy3v4t8/p20DiHUEjdxaafEiARlvVroRV4htRxun08l+j
6Im7cOO7z9kGQLSz/XboILx2U8Owus9SHnT5c61KXZqVmBbUfpj/XP30eVywJn5c
ckk/VE4GCAYZYaGkgRkjHcXi5QIJ/k6E3W6dueG+25T0GE7NY1ECmcdP0fN8qfxl
xMG7UIrwlAfWbm9En4siH5YNTBu8LnJpNZivenZbIA520YQiWp1QxfdWZHuwez8y
9LOhyibIKTFgIU5PUT9cYbGHvsBQYq5HSvmrFhGqM9+gqF9KfMpx3YLAXQxumM7F
BgnNcYQ19ByDw0vjALO/LdKCfj2BxqEs7c6O2kXvD8MQNmTLaqEGwDKYPuzojITp
Li2Ez5rdpSWYmIZSyMP+dUxntHapxR1xZcHKA6NifiUScbFJ+HVUmTdW3IWlnXuA
m+LkFjc4B64v6Db8De98gCYs/vqKwMo5NgzxxXVY/eZzCZZHqADXFM3rttQgPXA+
cx5ycwiIwvq1jcjeH5Z65PVkambgTKOphpVH6hV8OIvUtRa1nv4GiHtHbEOokkOX
VF3ZxanydqqjqqDffh+4tka3vDs6NTD3NnT0sc5vPbr81dZZ/piNaIGTGdHWjxAg
E6yNLBW6cDHX++IkDWutayAoZBt1sk3A7rNSfu0V5dmcAxqbJYMDhEyU74KzdB5B
qC3PE6j7qrH7g7I/8RaUssqUfs63zzuYl1ZIJZ70+dBVIQyVCKNlolIGM7m4l1+R
UQ47Y8+FyPpZF1KzIIn8gKkhTLtRkdTtjPS+Ce7r8qpJWLzSe56OTUkbzvWfhmlv
soUmG+Vxtyn9z74DFSitVKti9QAHNQvu9rv4dSw+CsS7R5GqgJcXD6T02XFPIW7I
kU9RQfmNpPkUANwxhVwMXZ569DyY26+UZUkkM1E2UBhB/jpIVEaDCXgsW33nK6dH
B6wLrH+e7GES9lTs7KQhSVKN0hd3VVZ9Jp+nWPnPiKJvhy82GimvbenTx26aZOpF
KHd0k/AIvqNbwKmJJECS31Re5gwsISi9T+xMQ1hGZy0NzDAyLwGIPb7zMFxtr+qO
FOZYFVTqCD1Xjkv8G1Y0Zc77xBD5P3j5THoaS9Cx5eX6QZ62/dWDy2z4LAQzamQz
BDZa8sBc5Ah8X+291OwQQxH1KIqbA7uPJ8LS1hIi23EnMy2KZgbIpN2i9euTw1Qy
rEN6HNmdrebPYAKYblkH6xXwv7T0ogk2/yhzTEZ0uzcym+n8K3/3FRZkAHtw6Efo
VxPNAfgznRd1k/sM03qw369uT2bcujxvzW0W2chdxGxBc3zrC3Ued1r5FKzlxpt7
vb5phLO8OO6zHSJolhGlyKpKQ49fv4Z/hfsPPpvm63Vf1IQ0X6ifUa5+QbWDl1XT
xUTpMnp+th/78Vr/BBDMnUsXPJOrqsFJjFjzhoHg6Kl+3GeKaBT+/wVlOE9j1Euj
Cn720/3iN/6uv+poofbIf610Omvqv2vP1QMt0mPS3+Qdoisw5GamlIlSmLXvJ9+g
UeC8C33iA4jY8TfiGGZgCfV6jSuf+Y+YHPQ/pFF93rSgRzsRT1ZNB5IUqoGA95DR
vSUnfUzlrcKHJmYEwLwApZhP0N7socks+mJEY9zbsg5qEvxpWZ4y/bmLFqOMEaFp
LMeAKEd/IKEOuXMe/cBLdQBos7nENL4ELh6JPupfM1PCd6V0TwOrzK2yYMBk4ufN
DZKvd1+fNWetVXYCUgb9uR0NHigXA8DMqiRhc1yGYNTL91M8dL0Bo5H1H0bSP3FR
OZXZo/4GiZlxjOoz1CnPM1PGIKAoY8JeuIQDr84W5DozvvGLyi+fksAqcjfi5cMS
T+m0GDNItcLmIuG4Mf22kK2LVIauiRCMhnZpNq+9pVuA++gw8gW6oFbqmtzpbOJS
gpW/lu+4c8LXOiGsIXPlSDBC/kNeA1bs3mhBEfkRMXOwbrhqNHM/mL1HUwBN68wg
iCadCbKwFaFTXUrpsZ8uQ+46TCxi4wRvUAz5fc7Zde9MCoBZoLp8UI/+XtWzHD9Z
cueDroqKYw+PRMbu0sFqVlNK3mU+SDl9xgoGSK7kxD//BBVLBG9iITmGIG819lof
dKXJcFavn5sK4CNLyCOrdcgOtqIznQ5MeNDUXDtshyfj3q5tep+36Hzb6yjRhbFv
KRRg59uPDfhCt7kFjuk49LqJkf9+56934fJqQsgTU0FkJLllEEQoLkZf+XGi7Hyy
638W3ReakOTp1EN1QC3kdiOfwk0TtMyUp/FrPDKl2upl7f1oLoC6mI3SwxO904hB
CZOp4CY1cIYH2oqAEGLN/y52fyxS0JNkjaDAE9IJ7IRPC8opwu4a//NAOhcfKOQF
p265a186ACXezD2uGODnW2K1RzsbUslSwS+hjYuJkd/+FfLPrkO2mHoVKCt8MHzw
gft+t9GmJ6NFcrsQdJNcRId7eownXPTu91Sr8mPARF2iNY+3+5PciQUUYgfVRBgB
a3wSZyeQbi75fzsHAr5MZ3kwk9ZICuIrxIUEtAoIMKOcWlmXxExUMHNvkMvRIqI7
mkQgYiBuZwn5cDijGTszRwYANJfc4V8+B6I5YPvOnnQ6DRtEmvaDE5FO3CAMIVhS
Qa/PCdyWuU4DEs6HENdjaIyfQ+5u6mNROBZeNfEBXXODerAf8++ZUp1hpjj+GT3e
TclfJpqHYG4XCnjxkSwdWx9eoR9iyfTc6QlvfVPQm63Mym9r6s2bJiQeGYKhZNUZ
EA0TdeNoilszGXGd03Wjg2icKR8CVSRXEzcdxYQg9zBH3+05bCC6fgf7nBHpUoTQ
356fdrzNDIjLraz+IdNwQyy2AzBfombHuoubKby3EcOwT0Ale7KIbGBGA/npwJee
pWFBRkkto7VFTsp42hufGKVL0FC6y3EYZ84dZi8StMWM1OnPAfZU7/Ro4NhRpNK+
FXdO/LQLSwEgdpTM90/F7ly2c5Cn7TQO6Oz+iQmXQarAoyli5UY3Kh95eJ0evOOF
ytRvqk5P7Q6D1fOxDr6UIStntL2kwVmPE5YZ7OGp6WKbuxDq1zG8jzyeFitwdAEu
iZ7Xtf8cHQZiRfk8sk4ZqhPdBjXGqp0/jSzbCpGRl6syIAPq4/NgqBkFoMmuek89
ppeFW+SNO29PblhR6iHBLft21BHGXYOGqImQVlH+6pVrL6MEDXOXBFuC1zWpAIHI
zU+4NF75bicCUWKh0qShnosDdtGlqKFvBcYS8gbF1ObTV42gOzJtW9VPSmgqtTI9
oMXZ7QPxAHSY2kKuzAdgxnSReObszGB7A8Qx0smW0cU2GRbDG2hOvgvT93cH3nRl
i+Uk5qShXnyJrJNQXjHIwL83BgjEajeNK0/WHC2WW1dJVh52SCbYMyr42NawKCJe
zP8IqXQNOGojIMzE4a76/DnhD8c2XOrRz70vOeIDXR/KbNfMuzRADYEHQZiCqTem
vpbDEK1qit1QEDiw4liKCCkLdjt3BTabtAD/3nzLhCCpXjxDwogQFtfCg4T7AUwA
/kX4MJMWbk6q0YIG/+8QKWw5Au67rScOTAxN6/MjsTNhmoD8W81p9m0U5GGQbhR3
ystesjwsUE9e4zapRqS2aVFw0beaUGraAyrR+WWVJ4sBRVGfq+/Zz2pLnBAr9CEp
ONdo1zMS8mshgh/4je1sw+KOxkZupdqcIDYmhz8tisieHgUFh/D2q9sR3qsKLxV8
2+Ish7yxHJsWaO7oTmWYM7IdEle6BUBIUksdkHivJ57I+SvA5hj4UPDYJewm/eKn
d+fN0fscmbt2fs8ObwkFirnWUIxOcgMFj8ST9NrNWk7QN3ESP3ohagEbDNIxPz8K
dBGLvGJ6mk2DujWNKPX/CvDY00eWYf0Yh0t8fzxPJu+T3eW7hWNY1fOY317cab2y
PFu0ZZW8wuRh8O9nfUFBGmNgFreC80tPapVVHCtzLcIteEFQ7ka4VRTXKAPG046i
LFBoNKNhIe3w9+PejGlSkdARHodL/F21+Pn4Mr1ZT1qlAAUJ8+gvJ+/NCycFCK0f
UjbA3IOfvYGG0Yv68ayHoLA9zQEG4ya9bq7ScRyPiHRfbg81xjBPrI4dsfPRXGuK
1SUYYix6CXJM80t1cdPrYjJdUQ3RYbD7SsZv+s3P5NFmpDbwVN0jtiOhAFYAM7K9
A6lSORC1uhQA8vEe5fiisai/Ad9pFuuQ7v22WtGAHWUd+sa2JL00BdY4SMBsm3/p
asEV1Fau5PGaHjPSMcurPGHyPZ99/5WSEJl8UwM76UyWp84eDRCEDf50x/Z35TKL
YXksPFWaX6W79v1smf5ESxZA3uzs1OVQjp+0qG0r69SV3G74v62KtHyzcgvghDJw
6at674TJOoaFC5c4P530KgW0itzAFJ2kMXCFDeM+upPB0XOd1hsumZZIBTdvP49Q
jzgmDVZu+km02TKg+Em3TDHsRHkUkvXnGRpJGKxYQlX+VoqkRiglh8Uu65oLhzZs
BySX9pSqiRiT7nDyLRGrUCVDHEzRUsPh1SqaBuKX2KA4inmdCSGkLQT+yl+G2ykL
DcghIYulkoDQxMOxmlP6/lLkxZDtqk28tpUVpr4Jd5guwL9jvbBTltZ1OpTHHCqD
06c5wGTSHnl3dJ1SFYbrmp5/QHPSHCFCccKJs5AFMTT9Q98I9qi+Kbr+oRW/OBd0
0fDhh/gx637ncP/DYyigXDp2xGK0CxoB008gwEGLwfESKMgPScpoKry8rnkDrWka
YarS2Gnq1XrZz0DEBrJFavYOpcorH4XKeq4VQB5FjdeLUjErxlAEErrlNJ1xGXSz
9U0npXnIJYtvt6fK3COcUX3QMJJ+C436tLdo/eNdEgjYwOtUl74VEj7KoyvCE0jC
0A0eL6c4fAqo3k/JQj8XWTA5a+YTI7x+8WSYPjchzcigeNDfEGhYIB702R8vbR5j
AA7St+DNGd+VDokC4S4NtgUwgYC0PlIfiEHQOF3yaIKG7/h2fgS6MOgqTNo4mapW
dN8d0uT8db1NHxVckVGeml+5dEGc3JwPT8kuRE3xesRkpEgYLcEOPhF6Bp7pWcYh
NB19MWZT0rrAKbJ9M5d9RnUAjeJbWsnbd4uOzvsKbvs3dphHkz5hENQC4LRFD/q/
9xHiEO2K+5IGNxyP80y+j/wa3FcpMLRb5XHmrttkZAaRImr23l7hciv8QUPqc83r
eWPeh4SDdFCWJ5fyzDwHfqjiQvIHu8lKq60pBFyC0J3eilYYlJItb1PU/cVO9IOp
Ar3u55tbzZCn0yHJxm1INS40CwOfbm0/esyBykWwBJTGbDYILHb9wUbYzsFV7U2i
8vxRGWVSXCi0ZsObWf6T760tsXeXqRR1iywS980UwZvXMyqClOtDXmK1nacD/siw
BDf2A4Vb3By/Y+z41tdC2pizssuFPUOlsNRzoly0dbvSRsIDKXvHfA6jBrBcEPd4
QEkvLCT9GKEJmLxTdsu6wyRT8TtyaUZPAFGYlHVW3skDaS+kXhQ6T4+Zb5+Z8mZt
/u1ZUgQSKvOsYRbFSewXXwA5YmTciB/8oig9lgJ57OgBpmAgZJvG2rAZl/AShqHD
7qytv/nuphAEZGYNZunRMUxI5wmIwQu8gUbvntqYBuL47P8CYZB+LYCrqa1kRLuj
rJxoy91IsU9VU8KiuBel02xClQYxR6uHZoCER9V3TyNECpJFWEHRMWbjcMsSYMyd
K/67tNGSG8R9KFgOB/27CYLJwEzfquJzffyTuECP2xRX87n/75rPTIVHUL5ojTtB
+x0eXtNiLhOWg26MpJ4wdR27xpqPSWREvgifa+OC6k5Ghu1Xq5OxV3qVShHWRbB8
t5abnMtFC9EfJXuLdcC7I6+XKjAc9MoJuPEmO6Qtw82V0cwK/EpQDUCvMkRcg2Qp
DQIuoaWp15M/KZvEC5f2kDElEzSJS7MTWdaXdE3mpRFqCHcWPzRA2QxRtbJCPaOe
uWCRcxGwHgPyJLI4+/fL443Hgcvw5F3yb4YSCIH88P5/oS+/HS3yPM/VOPtotIdv
2z+MC5VTysnxalF6R0OOvYFV7EbcFsLFTaC7mB9hQC6797+U5MDTMPfDhXsI3QnK
Wz+DAi3m54hovgpjxbyxG4Y464xdZfShGuKarLC+DfD0D0GO/yWukPlJoi0WSZ1U
P8cJjB6jkWzgvaeOSuVFG6N7221JH3kGCYzdvFBfrSyHloBYxvIiyAgiWBjauokP
y0GXo1bKhL/fFfT3is7d41gVsWhI3FEYCnXutin/wCvrDvZye8SqrPPOddtzqSIE
3ZYoHXuNm1ES+aF+V+a7iWrK3F6WXE2UWC5dcKWEUTDrK9+SlCXjUIldCVsY1peN
r2Bv2uJwIMcQaNcuCBFhZ/A4+gfiVMhpw+MgHT5Yh/HzAm4JkVnuhmhGjSncnISr
VaCFnn5KjUh7KFPS0lB1/TC+RVPXFSfip0cvJfFk2A+9a1Eb0jC4IyJ8ccbwJeRB
Dc6EueA6812cWyoOw+xxG2Z4bSGlT+yTvaMT2R8R5i+tl1ImfbxpAZnA+S3qVkfq
jy8+LGCOLcE658O90eCfsIXF8oOgtb8L5puafAgQ4/+smN2RJL2MuFwy7W/xXpri
SbscyshzbTq9Twp0zvbptoE06joYh4m5M6xkX52Iv6wd5UBNu+Pu9aKbnCUbb5xP
zKPpjPewuZtRJPzJVv3i0keYlbPSaOUmJt+XOh6rA6HFT+PpsQJ7tzKscU/x1FVK
meQBQjoIgu5BMXxeX0KYVPyPRM3kJJAAok0bZUVXgYCv8QBed7UzuO0EmUV+EQnE
xaodFmuWtRDoHtQCYtssufNlyIJZT7eSuS2c7y9EH8w0oY3bZFQUZDe8LHO8OzQR
iVZZvcUY1N9c57jmIstB6CXE7kRwMVUKU9+TocKOTCBK/qRrhL+ml3LjSqEnCqYs
Bs7uwGbqGPmhlp4CbYu5ijSftGQpZ5lUXbvYL9/VNSyAd3i7ZiX9HHXKfM+IB4Ht
LsgjOWo6T+szW1uzvVb4F5rSNroULTaKNTvWNiXNqH51N3VOKZ+xTvxdOTDOE/Vh
V2x9nfNeEs5Qqm7UapHbe7iz+6SX3tM6bPaHQ1tgL9p5k2tp+7dDRcYYbQxFS8GE
JIJ1mzCwknVOUQjDv0w9Vo0q0WiFqJfZdfNpweKOxkMLUHVgYDKQIg4yHxrV0RgS
qDRDO76wYERnUKA+SGDl5tBwEJyGygc/jHt0/ybfJeEToD1nRpObqUckM9U9EWNU
Biy2VAi3/t+tR4qJJ7VYSy6AeUNzj3Le+KQB/vXq/r2sjY6sKGO8mgTaRccp707Q
X0rG0h91o3EktCt5CGvlTEK5+q7vnahiwKtCiI372O6xxYOKAGnZ59Ogt4JZy5BW
mrsq8p/z+nJZPBPhv6XRJm6VhYmae1YBeFa6M8Yt8CZ1z9xaHRBykB08SaHoiCGj
2D3e1meq4tGIhH9YTxOERC87keeqSUAaRX2CBsUiJ2KxOx1ftSOaMmDFx9O9++oy
570lqRUuhuVmF2oF19Ggqtf5lCUdtGiLpohN7sowl1aVCqH5VM4rcqANYrTw1III
qLZsB9wYK7raKIhuYJbJtXtK/C1cGLsFxCr3DC1+dAQ2t5XXJY+Cpg1rJB+UIRrf
XDCQeYPYdUT/uSdQvGrd7j6FLCblVI8G6XZaKMtR9SElPAfqUlfNWcyXgSGK7ZfP
gMFxz9GLwOgt4VIPI2c/nKIMEXcL2obbpISicSJPHOdVMo7rtQX9UpyqLkgq6R1j
QL0HvMMoRGf6aXHUNpP6zUq2pE32PiLkRjzqm8CAbnCJSDFtNffIdI44ZTKQ/YhM
+jgXX6EFQ/WA8glkvb5rf/oaScmq8PP2cPnDD7/mYJFu/CY6QrPPzf8kqwFL4bdz
9RhckLtJsFpRPEIJ86duFFLs0AqT12zHpTqpImeOn6sGwPTQ/oylujwXffejpeTk
UQOckbomaNEJ/NRwScw2JZHUn+1+reSFdl08N0R/uVriB7oD/P7SULjIgAL1/SkS
naIwE5eIfaKl5D6e4iR1JAjCkPBnqBnTpS/ytjopyNWuBr5GbPvS+sU82rgnWsj5
73IZBiEB2QETDbBcOtNKGMD9eS3byLnrfRpTeIxDRREg5UAKPx+1f681LWrL4ZTu
JQJD5ZzmAFU4WOe2AwfTJnzM4s1yLLLRyRBFdQJGJhDZSX1Z1bQnRJT/2CniqH3/
+s2RGavr9++0n2fna6RvioHc0qDKPX9hC33ErLHOl5bisR4R1n0UvYFLty0d3e6E
bJWD8el4HzhNCGMySxDYNmgCYX6kyXcVBqdtqPDXIMvf+lbMB/J56apX5FKbJyvi
2URZFtcXNll0XY9xVJ1OUjmp0z2EYOaGy9DlingZSAnWWoSaZoKkwTkJ9EX1Tm58
p/fBq5jk9HHsaL8W9nP0IlIkVqyUP5mAAZKKRdCaKXBotkgJvgfpjCZO81ZlHdFS
pYwhLcdimL36JLIR3ly1yOj/3lBQjddZSd+6yhMl5SU3GoH4IunAua4YMEIXdKh3
yfoFQR7+J597nSjb6XK7hp1Dc6cdOH9oEpFRajqRtKbh0/2YhTwhhtPifR8CgmGe
74gOoKwhALm4EKqZf27yuxqvDacdzMXzwg4SbfUoAto6Ya2l0WKNxHJZMfZJPpWy
`pragma protect end_protected
