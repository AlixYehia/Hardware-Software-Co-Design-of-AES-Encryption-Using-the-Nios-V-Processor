// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
H7qLCDR1eE3K+wfysNFoNl91jbro2rBIlA/MjN6ksgijGMSoj4AoRvX66onEiZqlsj0YNy2cyTW1
TVOEXzJSaXYm5KBdx370OaOJod7O8kRqfgjVkXwLKqAYs5wlt9NRoRUBkYMbAr7btCePmuG9FBV0
lEm15Y4dFmDKUK3Ni8eLMk3jHzLIgdBipnO1XLToHEzhIFXxPTV+8CsqiccwCe6PYG/yIumCfmb8
OPlDRiG2vksliJabjfgEeZfABqAp7pq1014ItmOS386AKIe9EuE3+Vas+FoeWBX/Mq8DwloEBdj2
2vBjlilJEuOAZM6dirElIbSvQMJiiXlqS2yksA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14192)
r0xTYl14K1vO3luAob/ettndQXKCHUOtbgnHlNRKP6VUSZhOK1xj+T8vJsgzUdsI4D7Ad30oKE69
pOO6N4GHSRZbGSeun2WXZsD7HVi7WsRJdYTUeALCq1ZOJGX0663FS0gS3+GA0iluOU5vP8sSOZFx
TykID2fgtZvgkBvKp7UMuvRC6YfWuppW+hJtVtR+VzSYoFfC7QRbN3cMzUwJvwImF8g0FEPT3b8p
oERn47TxF3QtmMRK8MNN+2qlndvDxtbXwFayfCaMBfHoPMaP0X24owdYlUj5chmQdWJUYrT7OeGk
PZsUXhFKbTRyf/65m2hLSbYmOKSBMOV9Yb0o+H+mU+mUJZ6jfW3Q/cjCKJwp4ERK/8n52lOc6HTa
PhB6Q6p2IpFfVFVMwaG+cRIwTZnBPlnMd73litIIy9otKBigwDBc8ITTsOKozJ1YzANqm3i0+wPe
cSOeO4wKvrzBOERet9nZ7y2SF1Fex5ilTCgP/hZwLLYviXmuOO0MUFg5yEstw/OmRKP7GkBRFXyd
Au7K52pcFjO1HqYEWfpa267RMn/gZc8JCMvjH+NeCg1jiEfYba3UozQu1tWo66pGyJ4NNSmoP8ad
f0NJCJuKprBE/B2ceoCSxmWv+KTJhALfO+/y5e1GuJ0iVzUBn7LkwiBlMvCZNXvFtrKsotJQLndy
zShhVJ87gD9j3TgdA90d3RLDWWr3OU42Yn8huICrJW2yIokjX3TVcZfigKQMGyyKQ6qS21y1hqnk
32CbzxOhzPVLqcTGvqScExw0c8rBNR7eyKBKLiSaEIiDilvg1wRIJ9ph2hobUQill7X3Ar2abbku
W7zD0uQ2cDhmZMN6JmtIp8MXsNFCiqt9BNCicUD+z0LeNFf9cXkiWRFyUo4/FAsLS2B1LP7gNIvm
2hqt3IIT96Qh3ZQrdFDtgbMnZpUmUMZp2WMPjgEOpRWJyANcD1CHDeU6nImHiuUAEr5wPetTnM+K
zJgYug2UQJcA/ZFUqSUBvz2fhXwzMnbLfqmNgs/KjBPmQbWd9CI4yHqOGgL6yEXUKMYwKN9mlyJA
jYPIaTm2gAx8oKCe3BW+KVfdpLkZ3Oo3snXlKhDV9lJOlxpPHKHNuX/L8VQyQv4rb9Fz4xqT/nI+
cAjQdDCPuHw+n4IWcu5pK1Uv57KCyYwWJuKlknR6ViBdcz7lNsFilYo7r6/x9I1gID5MHGGs1Sn3
RHhDTfwCANpmE1oqSSb3syC5Z3+ihTmTxS4tQhTJ2CHyxcclI3X9PdDIeuoF9ybW29ADdeNnX6vH
SwoT4UNsesQswUT+rGdIyXNukDUnEI3HXIgNOB7FoUaCYEj+noQzm5+s9uFZAB9X6/E/4C6Gs+Tk
9gwr1oq69xbj1DMREnsotxJmtHqpOlnaeMoQ2Xl3uWCIdkzlPWyyWN48O4re4ZkfoTvo/U1+46Q+
uvJoSFBsyxOqRsHf8QOELo+WrYF7nDjBacdFC3V8wlEAOsYuYtGvcPlF4IOC8lrsB2/MzjSdscxp
HGn04+fPQPK8/luXvNMQ86qI4B8FnkIw6A2GaupBgLrvRpuid/7QVeq2uqmRg2CIDT6gvBE1dkYr
ErUPn+RpJrJVsVX+lEJzt92Ty3r3FdhbWMu0RgEBOaXc5gjezkgOw2ns/bPJUVM9FDYjF4k7u2c5
PXFVB3ewTSdBkUu1Jg/QRS7HTioUKRhOH1931v9z8V/q2Bz3wH3Ob9vRLOoZf9BOuxFHa0H7vYwx
3L8GDSDJT9GrB06QU1FrNo2T4ecn+H07wdREcy+9ny5++ly99znK7RlxXyc2tzPnzl0SwEtCUIpd
4JEFkhkPzp25fo4CJp4/VzLjbM+itpJgkw56sqW4D+BjaWqyY965wliTJZKuFhUvz78Q8vngLR1N
M88fL6xOGGx3gS3xnEm9mn1NqR8IhJrMjuKMukFUvKWuR+qi+VKe/Iaw2GVUiaOAq04B0Y9wrMYf
IqDEDTViO8kZDr6wqsyaxTXm5sFoPavtrUv43ODxAQqKnZVzA7TApP2aHFF+id6HbV6tYtPH1o39
oOPmSyzVfkZslX7Mjtpi8VKifzQNORrqdVSpIuHSV2YzramgKxu9ZnG39Ww9KZYlryRIgWSIMIr4
LZVrYUvKNL9DJ+kgs4xed4UpqYqRYD5OWfknuh7hpC86dj1MnAUg/G7iR2lXSDJBGkLzEzi9J5gs
8sJD0DTNf3iQJlP8iecQslgldCaRAqBHMFqIKurm/ZuGxZbzsQDzgoIgihEi43vu9uq+PEsKLL75
5S6YfzKAueB7wZKK+cckm2LUqbgSxY/02qUNx3fWW+hR+8FKKrsnutfw8WXbxsSQSKVFVS8Tle6w
1z/D2C4uI5IeteWzQwZO0HKyG9mXTUXNqvejUPu/kyS8afZeryW7unD/64rU5R3CLciqb3KqQ8tc
HQqwKzrK89qTvD7S1dQ7nuD3ue7GaHtIgJnAP1/w+NG98+iR54kjikPMdNk6V1V/QRP7AflElaKM
SNt2P1SJgVd86L2Q+l+Ijs8sSCr2pElE4yF2APAXcHar4G4BFszgUHvmtmxpqSG6kAi7tqwdkmwf
X4IJaHYVnY4MCpad9ala2X6tbSBcE3QoDwQ4LhSmZwJRkAUi79xl11guw+4kCqdIh0LPa4rWR6ey
bAS+6M7yr+iMnOkG7rwc1rfSlXs9z9awrMm1bs0I4y7HtF0PdVsL392XxM7PBzIhxEQL4rSN42ws
3yF4bmACVCo6mVBgcAFjtonynbgYDG50fq2qDBK8tEVd2/JBkhmrYVRdqMSSiZmlu0FKMMgRQDI+
21StltENV8kH+OsFtlQ6u2Ren88HPi1CMGJ9CeARs8engkV8JKD5qsSsyzL/rWtQ5jraz0+eepC+
Yd0OPfPli1N8bxvdLis/BjsBbCPYPn7S5qumfS0Xs4uIBh3I2bvSq3M6m7RmbQcW6K+UMUWCwZ6v
wQoj4SKfiy0FCFWe/8dxJAe+bGgOlCUNP9D1b3qO0Tb70S9yGyY7f0Mny79PODZN75Y0fdWgRhY5
y7uXgvb4XRZMwmpvDFShJGe7yIqHyMHI9WXDvlqDYc70e5kqbX0OaJ9mKLyEdLs7vMR5DoXHllP0
Ey2rNmXO9v6SE5gEuLber1le9QKxgzGQs3LpmZ1fmdbTXPBhIvhkpx/Gz/L63U9dtsMuiIkPbxdH
+Ehzrz6yb7+8b63NPuyaOcT1X7gsXm+YL5/9iwR5yXb8d0IctCJPYCOzBwK9XUAvlk/PzEw0vKry
lAjgh/WAeeZtu7Q2tzv1/vz17ey+g3g4P5iOBnoLjpUtKHHiSQeD+opnorz8aUuUw6Mfc4MrUGpd
VWYJuRV+VFtp8xoZ61O0WEFaoRH0gnP3MmGZsR/fjsRGPHE+e50wsWivs73ZIf1RblOS9uoGjL61
XnY7a1uVph9RP0CatJnFfAMn5MFlxwJG1Asw8jjvtmy3GatFopmjauHfyieL90s0Xkbyg9rKpRla
WiHI9YlZUnY4e75Ji4O4TSTsR6VooV9YxPA+G2SHehTOAYtq7NUVVG2byQBgVe5mddd7W20aDC+U
xi7I2NAZNl4C/dQpDv3Jm/d+rMTslApyJTZJ9tye0te452ccqhi4yf1POdeME6kIU3E8yZACT2De
xRoD6QcmD6Jb/Gh5CxTt3bO37LbMNJBWRoOG0Q/caiyXW8NWp0USLCl8x4REDkotmsQqBty0f9CH
cVdUKdp0uI8FEOk0Rjraucn1CZYGBr0kxXJpltRjQHINhtnAB6hr5d/Dx1dzj9y7bc4Wx6VSwUfV
vdMxlmPGSeKy92gtamiY5JRWZHq9wpYREVLb07jXnM7I3CGoYDprlvkagRgV7FvFwgMgWIIB/sNh
e6oZyw5Arn8LexmCMcbgiPZEBK5geQ6Ha/iXGQAugIIArKd4OdAptrHkRKyfT0I0sPDJ0D0y/MAm
OIiNrgktrAZ8K+haVtbWr1+0NUdg/kXH+ncE61T29OovF2V2ISy5ZbSNbHaIf2yVCgrSUTMDW4dV
TWC9gvnM7TMX6Bb9f0/ljP/OC12J/QKDxfBlVsHGzLbvQ68Bp06zUsy6lNy0gOQtxaMM/5XypvEb
+A6+t1h7JHfwF1YlW3/0RWbt16h0eMzi4b/Dfw55shZ4w5PEVUb6BMbIa0up3bIZTq2yCaOJCwmX
ad11/VCID4ITNqPSA5P+8AjMM42l2ueGtqO6UjaW/duit3Iv43/MsEuuDR6o9IN2UCIwsoSafXZP
cNF71AN09dIP5xyzdtvN5Ya0m2fnW3Z/RPHvL4HA93X6PEQUKze+swhwYi0sIVQS9r8eienjiYSi
3M94lKM17/DNbgPf3f/q8DKxw5hUrPX+0TDF5/NEcEbB/qgeso3lfZvXGZvdJifBB+Fm5dV+xYqL
c1NvG9AD1badbEojfT13THD68Lrmru9DQ1Xs8I8kQCQ4jZe2Br1dozZj2ONWQ3+fCNOJUmn5AQ4/
8u7tQs042uauGjM7BMFmg8YGV9jsnyLqaYR3EDbmvGLEAVNosIsMNtkK7QaTwr4kqJfbVB+Brvag
g/tl+/hjMaeXw76OtpY5D/MyJb+qFHezDZhcXMIXMn6ke616bttEnenBmhdV+L332++2s3Fm4vqn
LYqYaBVnw7N8hcpltWcvMjvADjECqAf0D1g9xQWceJGbtT09+QTUfKlnOhWUjzHCripJ0OaaZnez
wYOocLwC8XvFJ69jcdEhD633Wd2KCXi4QKTZATEtk1Eaml6fXy8xriehgehdxDXEriGsXtRVL9NC
GStrU3QNEIC3ESI68aWd7QYMKqQeTSRzuULDEhML0OpjHIcT1EPSwZ3eIkYlXPDjHoQelI+4JJk0
s6MHRiR2KetNcE5Hp14d4xhNEmfDKBSvi/VIwtuiSeGUw3uNd05nzjJawJ3TETRZJZfaRuRnTtzR
ptQMIYQ4ekpVGmHfR5ikQ8iAI6wfLKCrYneZve6q3NiQdtSmPYK+b6CzgZ6XFv5PfG17xMVuaDrt
Uts4+mRqdEIt/uNm3uQL9h6HBug95KLExlbnHm0gbfJ8vRVnszEme5B2HV2Ce/Lm5f0jAcBAu00+
pIMD75fWdfvBCIR3sJ3UfVh/c+VJCASHFT0zaaDss5J0sB1wl3LCnoawkFVcyYTEQ+GK16GT4trY
iPymw8ozhggp6FNkEmfZmzLT92KXbQAVhNTTQ6WlMNnentZyzJJMXbMIMntEJD3zGpPl/FH9KBgh
6+ls6SRt9A0f8R1NLStVTq26xc/J/jNXtKeFWh00roZtO9Jh6ajvTB+RUfh5vjQETLZTQ60jzamk
MesX9nUDnsvCY8FmH6TAmDOu1gj+aplc5hXNMN8c/SKWansCPu7W9F6JohipxVT07aLKlMZpIOg+
rCPCvLnOTT5cffZtIrSpoxO9Y1MCG4d0suUZjtQn+FMst0JmHHqESS5u1sOfH2v1vTB1AiyeWr+S
A2GZpFWmJocTcRbl1QESRuvJZVZS9xbUiZmh4CsLz789bo69U5guaaMq28auaLetP+WS75RBDe3x
jm/y8aFdDuLhnMM9vRIoj3iPBCnATMHZboygvje7ymM4fx68zzwOs1+s27dEeK7FCmgg1gNmOju6
/msowmVWNiYy4o5KqsggeQVWiv4Ca+BKz4xBFhm/jgb4zJhmd1qHEdElrBCzKXpf56+J6Y5+Pfzf
oXs8YBInQRVQrjrPZZNEf4ugGt5N/GdzHLZ21RAM43Iooe90piB1NgSZ7Wm0OYIB4CwVQVbUA/Wr
FA1wevTQPLIv0tqlhOZ5r88mmxQfVQhhLfSqzqBBHAj8Jhsk6KPekIdm9vMdgkRLg8eznCNOEAdU
MzYIm+q/hwYUcFxs95LkEsfHQJxXEh0sH9vEQ9EBdVeH5w/nYBRLAp9EH8BYHyBPUuK8vOiAeasm
GE/fZKOUgwdQjAUIKrW52EN26yZiqxwthxRIE3MMGIfXxYPyJPLzFxPLyyyyQCt7Qdu93QitTSu4
lr8rmgeTBwlXC3lkTYNeYcxLZZ++2a+X5p1T0JGJ3yIadkAFCq+Rwbkh3cY2kO5R7C0tA9Quzji8
8U5RTLoAV+uf6pIG/oSlNKmvpmLB1JsDrjdUDP3CpMamwiZ+fSLzURKsHm6d97iV+6hcDPqvbV1J
zL1SrR2wqW9T19875v3eJ/UWfqd8Vo7iT3Spwqo/TvFhmeQRkQx5WR+qgkDCkH5+gM+KhrtFQmhR
7u0UasxHnLYemSTrDV+fLSR+MWzpT+5Su9K++c5t6WpRXNz7W7gV38EBNXvXY73inHTu5m0+BkT+
zz8FhF1//o5NNqY+SSCwNFY9jtfTXnopYSgByU+UlNozhZTfXB97MRkCxgXsYbOlGRjcWO5mfpQR
+AlaPJDziDOPhCnWqiJRnjxgp51eMT3P5Cj6HpDTOqKDQayBVY+ufwTFLzpnBQDhza30Uz8tcfyr
Q2o9x9PuzSdt9vnR3jKCSnG169Rt1HUAnsTNbfIfIq3v7t6kMZugwaVnnqWEfBuIOWZ0fM9KxivK
vpuKXAmTgiLfcpan8gqSl5NZMxxohNGofPQE/Ksaaey+TMHiXhqhJjAUbAjwkfM5Wh+FF/VMiIoS
Ir4e0B+nyn5WXMG89zigO+ISyva+EcFUMl6YCbIEIyoTl1+7yP0zEIzRI6WEYphgwAuy8LSkF62d
qov7fte1kBCqbAbQc4aonb01mFVewbZK3tZSFvI6e/CM+H2dRI04uq7wYPc4p3ArK0iJe7hzYBqs
oxCcpy07wWp7/DbiWcSpvGs9fT/aD/kYCNDfnvLT0Jp/vjlHQw4a3IRnYvdg34PQlUOnlIc+GBWs
SguBnTfrzsH/Bna2v0nhkBcWs/4wTTQ3syhSsuF6NUB4xGeyUJ+pjPDw8VSYNMkAV/cVlxVNpans
BwuKOGtXU7l039zGunh80nOWCTBdd+F5ds+podcPBGukQjEuSbppaYTdzU0pXOgCG/7+Nk1TJg7A
vnp2v7nkNzhnpsCf4wlPpGF7B1ndSqBR1ON/ISyHV7XZSDWzfRvPnTdRxIMFT6bOGKssf1X5Ig64
JT4PmK/nIVMHuM+YnaYcI9INFEM8rZD3PTsP3ZM4X3x/US3rrBGiDKvYz6G8YMMLREfxdXNEGdiX
p8Np46nI0B0upN8cIWK3YlodInc/+uKmpQaJGu5kkIt1AyB2mmCKsdPfSAb0EC7f06ePwbQyx8S5
Yk6u+JPy+cK7L3OTDeO6QAySAqeg13d/Z+1QhImavC+Q+OD356SGhMlm8J4iiPZ6oq3xp+8CloG9
crRLihWLHv3vgyk+/JcrjXYNXTZp0f18aGhajl9bzLF+HOOO1PTacOrnSxdjFiPuPjEvU6fiYAZM
LOYRt6vB0/QqAvcou5rwofGRxK0TKhHdb9xnIGlwWmclLacWqk3rv/QJockhLVUwrqM3CqPEHXxO
yP03c6Dh8M7r+wIJYZ9SzUguvpd1vHY//d/3XZIP+SgutGPkLrcmoH6X1iLTGCumA8jPD2DGvTsE
mqQh81q1AR7stgJA6Aqsw//6wu6RE+kZjX2thtWZGOLM+yl0QFn9LDzmQRwBvvbSbjLiWYyEyTH2
6I/sBMGia/Tn6w4Vbe92nl6qqu4QlAcv8v0UbFbKmlAQtbEXWkeTjAYDBUOlWyVBfzFjpRM2IUfr
cHCaiP1Ljh9ySP17Poi0WxbcXHWRxq2zooZfgBkeHZog3PolfQd6m5CB4aSe19ZvqUmEXxjIXk07
XFU32ZIByt3MBsNk1UlWg8RKtvA063uMblK9eqUN2rR4m1tkhfojZESClYpds7hFxfoHUke1yVyA
l/O3uUmPrI9JMuwhVYxNSITZn6T3CX8Y6wyXYSUFFdM+i8bDTcY5ZyFeS3xcinscIezWJJ1f4QS2
g8+pKzHzMed2/SEDsebG0qivJGtgFxNReWwijU/OEJgCVRIdY5iijpOvmoUK04AH9bKpSO45JDqD
OLa6agsGnGIcZfhYZ0MQG/tdFAraYYqcGSDMncnsytG68ouA2HqOC2i39XXqgPsbevJ25dhtSO59
tzijTnn3sviYf2Pp9SJbnqe+EMOfCxl/qEo5jpA0bD/hPmMgmLduBih3L9+C1NGGWmiJuQcqQhaq
wmwyXY74VuTKEZ79JBAVstkx9VqLLCtD+JcFEggK/xUqsQYMLGiWRU7gWAGzYappV1CdHHEspX9n
ZNvCCmpUoyjyV+OUfExPw+UJ5D+897Jr9w/ZA/qZAlwzbiMLsgJVJRCFsw9/KZpxsIoVGAF7v6Pm
Siur+YFcwjc02yEHL5yaH/UtajfseVncFpV74iJbyDP92JAliRnC4PEYI3a17EWrThbQXaY/IuCu
eyoBxtac4zS2jWJi5pvGcNAteicScLl2f5owg4Q8VIONeRIc3zBYWtiJcV2sfyUVyyXnIaYIhf8i
NknvtgvcQ223ZtSJ3bQcsT0ZyewVZOX+W9j1o9X+JVDyT5vJBCeH22Yd639oc/gstVc3yxztIKwY
0fm59gyp91zjScyLywN4zSrz7l/DMvMe6/KrkaHJ2yTcHx+SJdK8hyvs3PKrbnZrjl2WMQfOUmWI
jcyLNjxRaO7drKtzbZ1sFUGmtA3px/jjlu/9fg7LEiOW++zK4wR/gqeTAFoUAowptMsBovB8OvQ4
+Byg9/wKLrL03KJQiM2QxpM2gU5ZVxax3EAgv8m5DSCS7bJPndF3SBQJtC2FQHZ3XV4OlY6nckIc
nmzPM/pHiS1SgdJp4KtjX+p3GVrODAiZB4Pbt++UydN8dbaIGlpZHHIVglapL7dJphf8epbozL0B
nLWfNVVkGxJQ1qRFYvxBd8ZtLhQwJKvYWrQgklpMaDizRS+skZ+jQl2kEAMPgYWlkmc9yZ4PYFkE
bgZDum/5R/wQlv4Vgallria69EF7MAdeB6RPrxvnxvn4rfAXTEs9O916Cf3Xm24Km2jQLdjNBxF8
vlkwnWwq/tYPyJR+rWQTAl/pGvyKhHpeJA1KgRkZ193eePPOK5OxiHhJsVMactbc1rhBDk1W4er5
Ssmt6lrm46fnGvQtVpR4+cfYexfnUXXoI6KQlj7n/S/JtaO629bpVqQPwFQeY6TWHtbUAal/aOGU
Z6VdaeZFmbgbJRl+XfcVaYEtv1fPb+uSzIR5i2ekME6Yqi6qOJlZoDGDQRS96leHosoLPbL+Only
+P5HKlVpYDL/AYzoaustSZcAo4tZWhlTqfPQQ7M4CdN9ZuVs1vEeRTe64xuK14NLZXzSdQsVOIPh
biCqTABoEe4YCzciGdPU1+85Auy5Asa7FASGKtsVmCD99jZyZcBCNtHnQCePRTzhUEvRGvLpGB0M
EzQRf4nuw5VwQDT9q7TXGTO9BxRTa1/8yF9OJdbyEloMGQQBtlhLIf6O/+MK2FeeIXZ0K7VpJ1U8
c4ZOT+5EIv69do1WHWTmGUpohgCeiZ/yhrLwJcvtM99c8EzmxmEp49X97c1mVwpJzJs4Fup7Rv9U
x33bNNhyp8dj2TE6YrccnQYmpGTcq1BeKXtbc8KLoMQyRuonxwfiQEwNOpP8WdjTdQxuwKFABMME
0YzrZeP8M7wWoAPWGYUngg+uU5FClMm9N3FY3orjyo4RZamQ/xxMhWfYOPwre9a+EkSd4IOsMd53
akoR79wGUaSHZ+s7T794WGjapINH8WNfhY/NYssoMupW5vTlPlqnu/Lfw3tUtHVHIHrpAkX2xyEI
HU/yzncmqzStePjOEGcbdrVTnOKnHsnu+lPnZfyU65A2+R3aVm17198A++40z+cYK80KcOqeTI2i
cbmUekrchzSGSfss2KYntVBaHljn2BepFHvroE1ITFZYaiCIN7O/zQ13VjbHy0KuXaFHmKyJo/in
Hjf+BtIkNNFsi2c+oKL5vuf4BX5EGUAuh08o5BenIdb2ql81vSk/yqF6GclClve0llzLoZqDJ4J1
zK+A5E0JoshjF/jzr+Z+yeJyprV71NFOOW8kTnFuVM/cnyeUeaGsxGxQSnan789FFbjMGc37IfEU
KHbI4ngfpSNXvsLPJUKTS/AIjbC1dttwHTQKwNIs3XavHwdGk7z7RyQbPnkVkrZ/68cV0iuGD3Ra
J4EMSsNXQ5crSzUgmCFN7V1DDvKesKVidIppXIkuTOmDw/3zTJglw6PVEdj+cweqlUDyxiTp8YU4
AXYMyebcIKL0KLITV4O2Yi7r5XdffS4dk66gaNRhyYxttLdAqIwZz4UEOrgJT3ueuHgYfh7W7+uZ
IzHHVX/n32MmS8P6iSSx6yCncJh9aL10i+O9UUiitBzdo4hzMXkTyec+dfjsrNZyf+1hKgPi3mAe
ZtxgsuVkckaTQyNrmk3/7DIgDZDxLjFIGtQNRHTi/AOxe1YeoDz3edeDnySsc6PPQVrpjOiWIfUd
uNosXIRsYCCOlT8/vsAwVby7uJk1wgN0fVyRuHxyvXGyaaJ7kNRuvwHLFNIH8mICQV4STJInB0yl
ohZDCygtorHswVScxgOqqsad7eIGzQuaOYeze8DObetPF7cEJL3jKypGWHnve/d0/GZkMGL7oqJV
wNPssL1KE8giea6XW/FPfD3KlVt31ZFmdr26NPnaB0l0X3m6lOHHZmFR7ZV55MPn5+xslubr3b/6
+OCe3StTmjFhcZfdYGGtv2ioG+XK4jcyCkjsqLNc+hW0WwTy2onLTB+TWd5drXAkYAjnL60VkfFw
jubwwTTR3sHQYE/o8mixB2HiUyGP/4TbR4/RDPir6cIabom5+wRHH2B5UqDzYLPDDS5IVHFFQpL0
9ViqbHJ9wqEu+f5tDfNU0VDxqK7RlxAGtNvEtp3JB92BZ/NzSJ9HoDP5HEGnObv6F2pGDclWkVxF
FLVmBTfw+PVMLAv3i2/kyWArBEKkfiEHn1/4xC0POTxBDxofM2bsIsmqd+/ZIZwkVzqs48LZUIBp
jKKe/AAAGYeuLPK09gi08L4MdQlBuTDydNjFvEHYKGoVH9kr3JveMEIoTqL/mZ74pvWPucleGDFN
bFwujy1XUbBb9Bji8TcCBELL4Ayg0ODGLnWeXaOxaVSfZpPxJ0ncjTcks0rm/Yv3IzfcanxdO0ZP
MQlGJezmNQCC2BxEa+KLv8B5IFWT5gCXuq1XwPj+MmrDQn6zrvq3WhLVrsBsV+7s/B8+eYkJ7n8x
zM5WUZo9XsSd6jWSnGZqM9he3mrUeFoYfYHDkkGXEg31AYCl2IPP7Hmnu3ttrDScw/yg9FQFS6KS
z/l0mD3d2hq0ry6CbXzzadCqb82yhA4ClvNL7l6NPPDtVCAKdBn08wkWQsmkJN4sEtHkF5A/YEKP
EyBCrfFYzbOg+UoRahJJAGLksiw1U9BXXiQ+qYDJpPiYIDzud8mcJxvimExcicShee5SPOuQgg9B
9dbWqNrCL9zoAy3H0QeUjEy2jZAShBXZa6hZ4q9V5NkgubYFENsmZwNSXs0Hle5103DqpRePR3yE
lHgk35Yr9oVbaL+0+UYumGwxFtjCIjjGZb5c9Ki26ttWDlIH8IvCOygPWVI5JqGE8H8ehNmprBmr
fgrw3LgHui9KGBrFOkQtR/sPongbWlqu0Ay3GueIVcUSfr3AC5H4sl2RN9nH4hZzH264+eE2gFH1
VK8MJ90rJrLMUfkGXm6UR1vuTfhFg0qyMtk3HotNreayy2F8OsOqXaSUHTYcJ6s4E6E8vIUai6ks
V5b3rUVd4pRgQ1fKXnJJhuydLcxfnbiBApBLRhTwY1uh6oiFYg1Q73cQ/uhsgzSZpPMH1Vi8+zU4
2qP1vM5IoiA53P9LCAbJgLeSpzONVRepZ94E3dsQqWcxJ4LyfQcF3ApuO0tCHbtamgUKfC2xaaXy
uD2JnagPhXfcGG+DmeYR6sykekkrlgcheweotvGxltZIeXIeVfg8AfJ8P/ZzHwDfRzntGHo8cPrO
P7zQpE77zDzkQUz9jg52tpOM2mNaSuqaeX+rSTkUwsglIiNn3zbnEjrB7x0prbMzmUNTIb0oRsgK
QgUpSL5GOv8pjBEZcKG6ur1jkzMnr9pOV8u6iq4r+ohBzvI6Q/L8pbXOGD3JxrXyOTMCsjpaj3fl
ByRWfPVIllGSHK8xHti/U/N+QKkZKAx5TMjrrSktAt6R17VNu/QfMnlE6clAWWehL932Wsv1WjXD
8gQNY3u+MwA3eswVBy6LZuQBdH95RPF2Y1ZwSNptiHrdVZyWdikSIal1uh2ZKMueYZJb/KKgupB6
AOB/U82TcKOTMjXrBHGaCAnXVyYlcS+UBbyUkezvnVXu040OViiNafJkimogY7i2MlaMCP4kUALb
YViU+yreQmJde09O0ZaPQNxAa6K4fThmOLF9L2WtCtEEsFs1tkBY9UDYLOH99bQxRKkS3IN7O0kv
LrsKwuZT1ktnh/Hmk29cD9i1c2FI5XBxQn+mwra/NORo2idE9qrASdYpJe7M4OpBHZEQmNGYxz6y
YsX4cimhXwnV0UMyFcKE4ZmcGedn82Xjrqips91yVjqshP5hqZ99wHPsyXibH3alL7ay4ByI7a/F
dx09sqakXbQMU104s65KBbrJYtdtWqCjbnrNFJaQ5JJWxrtox897miQ/nnJWS5ZmRYusALyqX/mp
VHTAWgetH0awfIuh2nOni/BVOXPMZ3YN/13XveRZkC2kHxSaNkNYJXxWp3vWGo0yEH1Kt9QkLXvf
mDD3dCrleFIoGAup2yQUqvu6dCvs6KjIQKo+SNnfgROZ6ywGP0TiNY68Vbr9wJBOmwhi/Fg8T3pb
7M7Hj0YZ+JW/3i/etV3Hg2BpmkrQOVQ+L5ZFFcD1eSnQ4EnrM+qnhzQ9fA6Ev9Bb2DJS40ljSMl7
m5yWoLoAgSnS12E8D3Jdu6FUsU5QoJ4bnXgAceprEa3o4k9pnE24+Z6uPRA7+ecUyEo7NK9A/amn
JOdlWFdhb1n4xNirdv/sq2vmgzZtUQ3+6q6HxLofAOqz5OuXcERHZhIBfmHYIFdCFk8nrTnNdane
VtYWrUr/HvQiMYSmZcVK9l2KDVRIqKxgIQBolSvxTqgn+Offe4jeVtNbgwea2xPOOIcevNVQavJL
GUKr9fzjKCb9+65iK1HsgCXMkGrDXqZpWOZaAGAOA7N3WIoB8uZT3EwN07ksteQIQ12LdL798PPD
E8ZAJLFgssdg45gy4nXYV+cfX3KVNTfdMrXadTQ02AyptJqqAJDmvTQ5yg3V75osOUQfZCwiePoM
JmpQJO5+rdXFBlF0wuZ5ImzonBqJyugEP/o3/RldYtqe9N6dZde2kbXQG/PfzSy3LgE8EyS7S7bj
TP4e7brA6U4c+OEHj+ptFY4WcclEVxgd6IoR/hZUputdxL53DaN3wpcHev5dxmZl32t6I2ebg3h4
HBnY1Y809Y4WOSXIiYwxL21JXhD6JlyF6lDn55OsjTfSzUVWTCvbTlEkaD0yVSd65aJRaxqxeY2D
01zhTzQMM6NfQCJuvdSPj1qVfBVcgjQKzl4w43vyuDO9B7Q9JO0VLnfGLFRO0Vwfvxzi6YfMsXSv
f2lnxSNpirg8KcEZ0mKdf396BPUV5geDAbUQ8dfMHoocxAT2KujR85HOK59Kmm3KZyk9ETlINhdG
z3uQJfp6KYZosyLXceuu6pyvZF7thoY5dB0zIDAQbV72c0TsLShNxItQG8hVc4FE+gMKutACDRTz
F5R/gXfCXQqWSWHgdBJv0wy8clUv/Aek77wkqCDfs1PwCHz++xbidQ118gvU47el8yosmW7Q1dd6
Ariz8oOf/UQTs5GBzd+iZdd8F7LRk4CsxmqTZ2/v21WYNd7kg3cWJRYlwiDINOGRHT0+fQuJhqdO
UgAjLDkMLnIO1GYpejdSNyidocAL3BUcUokMTUwkwoxYmX2hH2E3drsqqBnYYnRM4d+olerncG7C
NIP10K4AV17WFwVNjKk0tWHKbUuq2RLyUI0KdhfTSmq0BrA59ymkUnPuR6YFVga9U2f4m7k1aHXq
qo1JZ8KObi8ALKBPYHTf3bLdM4/FIvt6WhW92ehYBgt7Aztle5pYia5QMXQwo04dOJPrB1AP/ODV
J0o0urfL5/ki8HykVVZftbccFeyfEAUL7guK3Iw8uNE4sYB2kb50xB9n2jHMbY/PIZOaIq1xWVfG
ILWx1sdfMvHr5e5vw2UpqmD82DliW3sacDIEzhDK4ZfjZkg9ZXBKN2tO9Kz+ftyhHaYUjolCSkXl
mD5BRbxJDI9IqVFwas5yPDnlDRiFhYc+MCT9mJzuKHynDSlGr1tDxcTbam4UgPnJWwyhdH41bS/h
ymAMTWF5XScfIeeRynye5e0Mqo18Dvbzzmw3LY2tGGej78JdKaERip8z3pugnQ+xRHoLh15w40AR
9UVTBRj449b/mpV/aBOa6Z4uaoT4iimrwsBoHCEFWzdYKFdaPy8+TKSAyr3aYqKJTAIQt8217mgx
ksATKEbgM73Z8/HfcP9oGRUprFdkZIwwZ/qfhNQZv7qdtbpn6WAn4+CqDsKYGIXEWiVqkyuzfqp2
RBvqqiMt0x6rUd1pgWWA4bkl99UBeQIxQbb5R7p0xIYiM5m/mF60jdaZId90bQAVdlq/rauYg/nQ
kQlohWbfmpS+J1hJF/N+DUkpD2dXaXaOTUGYPD25PpbqpsdRNmgLKIFXJI+KicNpufHyGhvS6ThF
K3fCxyY3mQ+cMQOgPr8FO6AmI/kGpAbQB4xJZ5mN0VYl8AHxV+u+dEbSaSoHakAKtPJHkZY/Mqo7
YGRbJGxmbDGdrMkWS4hPmMTgpfkUEfC2CZlm0no4rz7EEJ8lS18SbtDlyKQL3VPjh/CzxvhhBdZ1
kayJjQoQ2TU7lwaXAlyOlY8oqsul0jS+B6O93Rsx3acAAg+DW3mHlttd7c4rs63G2B5OuQNZ0MNP
denGV5pwZFLvLmcGkedPNSjvPWiTrUwPWGGj8cArSCZXbA0YKATKeDYfjWHCPtsEmvJD7IH2ILC/
y9eKZfg9FY7k77Qs23oyvJ3ChjT5xVK8T0xfrgujQJViVjBvZ9No90P8gIkajhl0JOn8jcuhPJt5
9QEqIClP1+gybcuqNP7ipCku9Ztexm3nmj0Gtw6CCNEUWOi76B9LgnElEHtoMe4eaitNmVDlYoUk
N7Uyhz4GH3RIWXh5Qxqk2Y1IjAhhGfADg9Z7zsOYqgxLHmFNaKYp0Om4notiVfsOqFJI532YcZAB
Yf7cj/fQ8R/OKPD9HlqD1x0DMM3f7DehqyfCgKuh4VCwmxklaLLZVWyy77kUHhUv/oUkVa1WFrG8
ehNiDPysJfg2V1z25PPCTp9O2CMRG6rqS0Ei9355IGtjJLUeX3Z8VW0Wd/s8fOKV0eov+PHugPTd
ffwxK1aInFt/G4wpIXK8Oj8rQI8wpqSEPOK4tHjbx7fVovQ2WpP3jXNjOk4RB1MtiBt8PsLhtx0L
laIRPNCGH/rPS+r15xwM5UQqiOZnuWFoCo/gT6t/vPFe+sQO6/1mSdtu/+fdIsnLEkuzrsZCQnCk
uvYikGrFVEsawsylsOgR2qAHmzhrf3W1Ne8/POH5Y52wFld8acONPJ85yUsYy1QBGZ82G5flJg7o
fSZAET8ks/fqithC+rJ9ctWyOvvKVzbcpbGLTZ/me7BR7JZY9sY4EXgwc8kBIVNoX2DanC/jQNhv
UwK20D6QyHRHjQbEQpDaDHCzW0K3PTHLROayex6kDlvofqPOWFtONinCD1mlvK8GReJnV8wXMfUB
c/ctz0FnUCMcuMnpWWz0mc/INUiMvtJIQbU4MJSZ764n36TMTfSGS1uuQsHeCu9dzgt25W/URt+T
ksqGM5NXbaSnJIjDFsjZpEBxx0TTGFKiStB38PjVAtt4Fg4W1aXh23bPU4R20VoK5AmqOrfRKU4+
/jB5gxzJsPrM7j25EczoyVv6S1Q9dNleK1JhlX0mZzuG6KSpbW0i9V8zPbqd5pHOgZ2wYZHqIvCi
orR8XcvsJ9jghoum28d95KHuJQnLYB7MdMnU+Kz4F9x7yWJF8rncBTz8/u3sm39KHoC/SRmCyMUu
SzWQY8Tq39e6q2vLNckCY2SjH9m0EJOinfJd8MwP5Z46rRgOPnJmD9NltXgRxjeFoRKIUEhHrT0H
U1LmcA6CKrAxoFt6HhJyK8oIvf3LtgsgvIGOTHsm9HA4aA/uNhUlSLfrrDugeXc+XmlZy4J8oYDj
9C6qqiKBUIT4fQZwNUm3VHSg64zL85Yn4J+36SUfAoLhrI2kkcRCF8rj7E4DWHZWUyg6kE8mQWWm
MSnwLeRYZwYxfzW5z86jbC1YZVj2PcUW42Js032+i+zkdhsu1eaINPG5Kk/Sz1mqBCn/sZBFDkXv
UIiQukArrXcLVObMqGougk5kZmjEZQiIwk2R9iN4A9mDIyf3Y5RtkF+v6itdfxiI+lA2bNrcPppD
SvBAy9qQnn//mfLwFPBMesKtbbatZstOdskHQnht8tum/n4h/ZOU4MEwGFC4VvvqiARWAzXNQeWP
cq4xqGYzowyGrmZ7yCbvZR6cZqIa3mOvXaGHXZc8RIuM8GNqzixTh2AmKVE00bKerDKthhoq/ChU
W8SHgYEm3nPnKBM/ht7/x33+zT7mWMG5fFjpWpqpSJHdN47ydsMrke1BzhD4AHgJDlPTv4JkgMDJ
J6v2dnL2SfvpzULva6ki++tdoXpnz/DQm/i01gJkycUih/DcmlfWUrdGjwwHsDtvz/OZ9ai7UtCm
KieblhWzsKV7vzMHTugLKHE/qQOJ3PhE7TY3EXMIebed+k43NRNFHXGaVZUcmOOnUPWXnUQnqA9R
aX3r5dTZsU6dDIB7HvVaeH1clsuhWKaF1jWSgh4sjNbPXEmXF0VZjuwfdtXwy/gZyYw0bVz2xj0T
FoKm15HsaJY7ftLhQ8uaThLz54qU5y57eaoD3ct7hQn/Y2HzACtnIzK3N4exMHwwHSzMqn0+Cq44
INT1DXw2pLOjGtjKZUjLNICkuYCzbVJq9xLEtVGgecF44GnAqVEf2+/up4aD5NKbdAY5pfdANnlj
XMqPGwnY9gwLxxxv0rbpewzWb1B9tbkZ3vLsR67pu0rJkQcKctsAc+E55km4HkuGD/15XFh59C5Y
kDhV6lTvqAkYk8JcsgKWp7Ucq+eP6U1rsuGbxHR1ykJVBYqtBW1Q5e9aSMlH4KRfx+0hcdiJtLLg
Uozo9nX8YYlX4kvQ0f3MBMp/lpjFWomWSOQSyvjNxzRGUxNURi/tQ2IpIv0kMfPH12ADb8QGuInI
g7zqkJ/bVq57m92/Il+YVnkgXjaAIYl02fUspLqDZlQzEKOIjkaVmiKFWwIIkaG3jkHn2xb8mLSx
un42wXbIIh6emR0eq5kswOMgTWcNj4AiXR+EcXEKhT5DZ6NPJWELFzxzz0AOChZn27Zn8Tt2WrVK
M2SQcP4FZZobpf2buf0RwR2iK6UN7ByrI/BwFW5Bz6EMrup1LlLZDDOBPNBZKuK0sHDwe7b8Fvp3
IjY6aiFIiQF4GoRzi/4dDqdV7ohTFItm6P9yKbLL6KX8UyaCR+wr0aOkmiYP2f4WQTES47XTLyvf
7UtRuRSlaZj721pMAwAIGMRs/O2iRJ5ANdzG6PhVtcsqQGFUjps5+VFA9uZ5HxNomVh2nR5pHcr6
a1f6BFKgBFG0W3WA6vHci6Lw+aRbpO3k/PtPcjtjDiTW8MUdhJGWj8CQiRgGuUwcHR5aX7bGhkuY
BLksYyfsTYPFY+mai3P24bifvLxsCuP5nu+NM41sMcWxG+Sh6/JJ6lqU5M7jaqUnSdRa7SuM9cc9
s8UbXpTcFe8fngwds3l3965whxouZW0m/l6er/zEjW5EaTOiTk4GKCk+eGGVt4kpPn9pG/LaVG0m
r80mXRlKykSj2UUXUCM8cSY4L7sw0MQ6oeLiqzSuW3/9YFSuEVoA8d7k5eTPBwqH1AsdSDLpbCjQ
917yUUCw6NvqSbwu2tsFpVB084y48G+CtMudHHmDdi47Chnk3brmW5XvG5pPVuyL0pMm03wJJpOB
vCooLKjP4GyGIhiGYODHOhePsi479pboQSFtPBvbKYgkKOrWaPGPSWdetMeVTjASsx4ADe15GZHV
zS8/tunKXfsxeEL/GgXpoLtrhGSLen2uRtuETOlxEIXaZTuhnsUtm0Ue55Halpp3dCeN/Je1vpiY
UDGgXoa8KgSI4yhMbPJRFhmEAl722njKubJ1gHPUx5L1DxC06wJhgWAkZuyOfZPQl1GMwORIs2nn
1LdelSNzDX2go/+YK6S0w2DwfrtsKtv5ouZ1V6yeqDjEqc5NUb7tbvhKCn4pLYzqkYfT+4EHpj7r
WEjxSjEJsGDk/MSGWnBe8BrDuc7BWclDUu81Z1QkDtf5fcFxy7PK3o44BeldICNowshyInMvGWH1
XBosQnpa14w12pjyhllghR+B1AYnkCGWY47wS0Do/h7dSzd2T43BV26kE9vmDH5aRpUm3b5N9eOT
9md5gmWlwRqkZTsL/VKAqzCNgK14PxVglQYs7N1XmaVlTNpoW7cbHZlTXdHuG55eCU7ntBdeAYuz
ff8m/ZWAHopol1ODAPqe0gDc+nBYNrsLHQH1N4kSjIMXj7M04gT0NBcuNZ66K6KvW8lqCi9ExviH
KFqpSFBNYNk6a8dlTm1A7x1BiGnVxiZF2WxShoikdpgWNjrGo6MJ1qZBMGmb1M2ttrAhG2XEjnYz
+Xj67bu4/qWpI27jCGgEK7neNmcwCZByS+71oT+YDg8ybIXjVItHebrzoRWVi+igzm7Pv8M60i2S
lrxQqu9wIH/E13f8mEiXIggnVzueKLVNs9qckRkKc2nFNn3ryRwWdmOGUAuQyBK+gbWJ+Aj/uQ0k
XRhWPgKks+2MmtubHHD9/RJ+XnPTdG/TbcAEY9s5q4T9wHkvIiFoi60oYagz7LxEhQS/1dAq3d8=
`pragma protect end_protected
