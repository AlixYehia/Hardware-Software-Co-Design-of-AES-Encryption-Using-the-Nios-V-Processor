// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
zkG8oisrwd973NRkWy7sw749YaL2ORzkzH4avW6hk6UQs8LGeQabh6bST3q4cPIhMfCMQ7zm1qCO
JA/AdKQoaJtdDI92c8SWFiv2fTJxQzrbbMji9+yc0gt+Si5tKRvjNg7gZvb+rYGArxWB5jLhik/y
FgbY6i3DdjGzWFhYK43GAFCzpZWBPhVbFPyyLO4nRMPI7dBOTKZ89xBmzQ8njFTl4RPB3y6R02oq
W5ZD4JXVC9QBVRN6qi1g3mw7suvkZNtAW7vuqP/vuT1L5WXnDtkEnE6IxpXPT4RSHY1APmVuwK7g
e5xllErtr1kLz4nngDcY5C0JlPLTs81QfhY4EA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 49984)
scqjrsd9tnhGP4204xPns7WA9l4+MmTwKUEAea56ZYuR7PHWbS/W0Qgw2AGIU29gMRCscRn02tgo
ul6pYDM76h+hD/Xxw3NICOrcG/+PsLb3zj03QLDbWaO+W5eWCr1ow0Rezvc1hUcZdUV2FkK+EDqN
3+MxF2Qq0cbFvhUghyud0X4zwenBdcw74bbUpR+1OcGJNz1ptwLKe7u/K6ezhlCZlh+82J3k4FHT
vQB4fHM3MayA6tgyymz1BPx9EchsVdENPoP5RNf3RH6StKd/0OoGlSNORE+RPNq1jfLxU1EK9VpA
6iHEmNuCe22wghoaEGwNOQAHvinbOK+PISdACBietg7ne7tBNZgtuEJ7DK4MqEY8rqVj4qz+vejP
syZAL5mEOFE4fgJknDHOzSQgOGdAcoYa4SSvgiClFc5E8OkheZow1bqcSg31K6fa9xocbiDRy7Ho
yqJU2bb8FewaVycBtc0xppwXsHXb+GCVKOuenxztxVmFmNQbWwTyETqTfS6BRybrIMQQm0R7mD9Y
IJZY6DMy92QQAqqsu2zAV1d4fdQojBGQzWdp3QRc7YvqNmd+N7VRyPKYBknVw+mFGc5X4VBtsp5y
QJ7ooHI2LFQRzJ1OANShg8HH2+aKQBjeOOWfmOa/A3OSDbbNny2T2LyobSWzQGZzpHAQhy93jjvb
+1wYvYjx8jG4cMq8TOVDel2BHiNriZna6AaO43IEWzZeluY3Adbdc6wC/uRWQOPDnH3KDVp/oP81
7J+B84Rrpo9ctTmdqiIX8/6xbYaPDWYNMMBEMRuQTHTD5qowp5JsQnkHagoQdvkmujvZYDGBUnY1
2aGmawSQPZbH62URY5WMPFMbX1cVV+i9Zk6bjSbQJXm/R9g6xKtaHUNbbIZtj8ziVXCFYCQKHdro
Q7SUVJtWReY81GXsPJ5jUCjNl1VJMaWUapcI+Q34sk7QJ9BNETQiveaZt5uuswnOHQ+v1Ys2x7/F
sXEMjIdE5ykrnjCV8gvj5eRzRY5Wxc7jBVDn28X0ToorIedXosxEuY8r4tNu59PcbJG3O1Hs53mX
XZ33WbbBTjLxYaSTOMaWM6NN3zM0wtmkKOY4S2zgZG1XS0tyNp4hZNUd58nepA43/s/qSPMItyRq
CWlbWbiaZNLmKqZ7AVdpwfNvir6C2uHXtlSSI4s2i8c0uHEvSjH2ZvtE3KYs9LKmZMu4Yt1L3mv7
V/nXKvfbZwdI2T1d3BCShLoGBB388nkekQl4J1iK0V+ludjGuVXMWn6hdRTQttGqTXzg7L2qamIw
3ABkK4BI3v63xCXktwOC3mJzzujdj3kn4ecqHotf9Wd4bcuaO3xGyc1tIuaoTggRx4GDuZOSXyhS
cYEMXpvRs9Pk8ExDJEkBTdQuErFZhHZfwGnLEJ7XrlaXyOb4ZDgU5d7gSVhV5MnoTvTl5frZXXd0
qVOG/whrGS6qzRbDI519OVj8wYBgXePlsf1s0LumYwqT+8xPcbq7P8SkQyp1WiV/GOLuLMjaZ14w
jFyEfKF7f1bENXv00W6zxc3uSIohnrutxbJ5mgfxbFwemJwJjXLQiCAlGwREJZskyzhxjB+mIbLH
qOcG98iUuM7pHc0upyyHAVrlrH1jggfASxkthISuWcf/mtqlkmSsL5F1zYLHC5X6kaYfZ713FVHo
UTt2hA7iX7e+FJU+CuInRTLSuL/ew+OLxCskfRosCVGKv4QCBM9TttqPsoWulZxhnRLiG7fmpY85
AOmfYHlTX7z+De9rcNYOZQCoXQVNmNolfCUkZ5yDdZw0wL5BUvFmomqa59SWqyANp61UQbmhgkE/
3iHVmRG8IjqhpF0WfvdbHI/B6LBwZsmx7WljfJ9YNEdtZ6DsyqXmn88hH0VrlMEzxqNkT+Sz5B6i
zsC/euj4R2AgQqqt4TkwSxyQtE4q3y6KumYo84bv8pZsPZlgJJPkfU44orMLgZH+7n/shPh2FLvZ
EHmrLdnzTr+JE9A+iY508u75yJoq1g1v+HVXJrCigKYTzJSK0OfEJBmNbPL3bnklGERlhqWQrZM6
Mm6Em0ziQX7PXMeoj5upWyP7NeLM0oBjMv/q+h4zPhpRbjf6HKAW/3ZES5hOGLK7ENTR8Y1BG0Ny
fEk66wBKIr9UMlgUuMerTx+JQceAT2dZ9qpK30Qx8qp/sZBKhXL/+19LbLJ2Q1s83DC0vdLRjkI7
jvsZmd+kOyBQlRmLdAYyFBxlb9imi+qp3wMQA8NszNr5y9Ss/NqCXUrT3Ar64S0GL4Hb4ayhirR1
q3BwAxBKpbjqEikrhz2ELeFE3p6w0AXvlXuZQSomQ7fuf/E/yxBfET45Kf8i1hTwx0quOaJWG/26
TJIm+i4ZsLYzYT74oqjy0qsqsGvllR1XJC38cD3C5mYr2aQfal6EJ3UfmQTuNdBGkfUfvG5VN1c/
xhjpMSn1M1jwqXNQgJnwA5QUwAhaWjVPFqsey9ED1gLGcrwI+Zrq82M/lUKNpUlUip++Un6GNnCt
glTFAhLV8FYkNrZD5jmw77R2M2YALb236rdJ7VwOIJ139UYtNSN/TY1n1HV0R1fWGpImINK20Xu9
kUbIM0j7Q1gffVetI72AnoVG+KXeY3/5hvmLhAyIqB0Rp81AhnV9r/2xjm+ms/9f/pHEy+YwltuN
B2mf87o21ofxfKmVrHfeyXNasU4pmX6cDneHQQdQ0agSviYasP+1PX1LGWF1pi7CeBjxH7E3jYe2
SfG3dqbS3I/GvVZqsGCKvO9f+0Fy7z/eWa5XfVxh1uvif3FMcgrnUbDX+UtQRuzaxPTEsSV6Z6xS
DRd+7oNP4jyvXeLPWN43O4tWFlokxnHnvrdl8TmNWpgiJQw6kARLoylgih7Ky9dDTKQxLm0K0uXq
aGr53RDKslC2BidG0jAa611AmzJxHzmQ+vYv/zlnykMwQi081Mgu3wvkJexYXE/WCzkA1Jto0ElW
j+9bZmq0gQOIvTDgWzF4dilohCcgNBZgNW1Xu6KfWovZDVBfz2WcQb0hjBg7shAbXcdvxq+1IclC
xYvfUXNF3p6L70+YglC0f7NooKUwfA3g7Lu/M0V01+2AN/s+PF6kJ0CSt+TNGUtJ8v97lxgOxqFY
v9r8yWVOo1Sdr1/ytXCoYXUi/LdyDufWdwcgwIA2cGUNIYtJ/HDavX1i9oQpHlZxShBPJhNnvdN5
AE/vVjAmi/4RbnLrchyL8/a4ylfI0uoEawQBRbJYUigHDIRNV/uEFtIf17F1/8M1RJTzLMCTa+gq
1VEjbZoJMNQlok8P1CBKlqolD/R+qbuFXtbCf7gP+k6xtIzshB/kGMO5nhuVk39IjcgkSEpJ3C/S
vqCcAUqNgmHxccpzn1MFqCvie760YV2cmHp6sAmSHBRmFPw6lIW75qrl8CS4QtuUAhs3ki/6c4UV
LbfCsg6TR/oEqWL2YUiEk7VVQ0lTHzaVaNii0S/ibBLcUjGSSI/XDuueH3yCX0IwGLiwU08k4AAk
O7iBeD7Vb5IgUNHBIECkP0QcDOswah4yN6bHoQIh6Yc1Q/t0Gv6ScG43eOjVxhTI8NPg81CKm+72
JzKx9NFYPDzGGmjYj6TjNGWYCdBkcHYEHk49NkUQz2UuWv42VAopkuuGBh/RiqKRmnPsl0H+hZ54
JIRr4Cq3z4WLl0uO6SV2ZzRJsn0xBXAHOUJK5JAD3wz53i3sx+fgYsBkr280WV0HJRgRDinC1da5
MTsV7fJdcz5isDCj5QZPcmYnJW38Tyfzzh1SjMQeRaVjD64aNyZdfmUxWZRac1J/P53MW9VGrFKC
FrTvas3EnaRd6wmHd8Yq2LL8F8ceK1961uT7TSizz0bsp8B8Z2DXocCy0017oMyGPstdpAcJBRkg
i+RRAPu/simbA/YMcv/9KLXgJ5MRxygTWi5ZIIAFB1Ek7ZEajaLO0yUS8AsDg8FQR3ZD45ri5xI8
Tp/9W2hzCpKU4EBR/eU1rv9BQIRY/Re2ALAwVirQUC06ix2T49BvpHDrRyy4TyL3gqgexPm4ssLz
fo5ii4AFs+r66GUDLsVkq/9T5KDMCUDPhprmEa/2C1SafI+lW2/YrlmawbJeGFqdLkvrQBNbuC/+
Jw/gywY29ixJP+XaXrRkApo7JLM71GXbSaMp2fg6ezR0rG3mF1xV8UgEzm6Bte9bltW4UOZMY+14
/9qR+dq9T29anInsACq+fwfHDQouYOMGSi9CfuIHXyz4dhJsYN/zUWv02buiWAUziGu7KCWsQXnx
H0CyWw77bM9qR7XyLAGEc9Ef48CSMPj5Y5KLfTL5VjpwIgtfXWHcwLbX4efxXzug4n6H3tjOzLk/
+S+xCAznJV3jC7e5LY/sVc0MRUPOnmatVJHtMkeud27BgY8ym9WGRrT0++PJ5okWZU5YEejnWsT6
drhVSp66z0+3UVTAOLzuPk/hvdKEkMvg56/YNYlABsdWUo7YJD+kNoMis8dmZFVHNXEWG/0+gaIs
NjcDu3KIuIWc1EsMo4hCbuxgioAFsiSQnWHSisMG1DaCUutiDyPhg7GMqLSoSmvhXcD9bi+ORUTK
04ktF4ADUKGJCpXOyJRjZt6kpv1nAEGKPXDXamxOZqWN2RgSNFChpuldH8704DhRBPbdaORRH/50
Yitc+mxUJXqKVwawCkhBn21XoY/SmuuBJYZ36PsbB7ZglpgEgqv8FA4LALmk6mniPa1FYZl9TZfD
ak5M7BpsvASAEX6Px1ZDjMILu8bc5zCuveDfQGhX9rYANxRIWgrIox4o0ev3vYaZuR2vksu4rWZ+
LY4EJ/X6m42WjLmth0xCZ1aeUxaM1J/fPex1599wBtEjpJxECXj5EFCr4UhaB7fFhKy1rJNmk4Ld
E3cXpYuzrxHmVbVSfDQGtWZgZrmqHnZODCMujt3HjieU1gyr8O7DhhX5RGGNEB11APc3Cq18YFFP
yj9TKAzYVDMzQ8GMH1skv8JYxNuN/DiZUReQlZlIOHj+g8vhRzVSXrQfi+DS9CLOqPqUTp0seKju
jXTWfYOqV5xrBe8NBtJyWS+nWhXBB5u99ZdVszaPaAIiY8mSQFdXKtmAGHgc+RHzoY0ufosLJsG6
zTW7JRS9xDSH+ypGkfkKD01vkLC11nCYEP5ie/jcVTfgoPrWeU27ltjUAxvOoTdlDqT/DZ+paFgI
X0v9zB0/CZ66p8R0aY6zklntEJFnMB+i4AslHt2T8AiAZ1rMCpyR8hET/JaodW9DqxuazO0cFo2/
nenhNXDyj44SFN2x6SADiC6l8h24Ca68/lbe6nHUXMQCFzdNwgJr31VvsvlriYYKUJZarrpf9GGS
9JZiqLr+z7hodNzx8p72v0Bc9si3peA46CDRurYHmTXQQQSR1gInQ/VWyCx6+rGeJ5cqfYq87E3c
uGJe+ZlI41UVqeizFqt1I9+6DkLsM8DodWyCRoYbDsU2uYFC2ReBdunDUHAtig7zzvHtZ47GdwhE
xSUJaHeaJcqzCGwJXHOLKozFK2Ch4aFapmGjy6Bo6kAQHlWhpPLclzImn6V8FHl49IJBJd3pZGRT
g/3Dag9Vj8FEAddgeSY6Y+0r9TxAHgs0AARf/3vNe0Ex2J6IrKm3c/EipnBagvSv+pDe5aBSeGOl
eHzhcmzdCeN0+t4Z/zwcmnLQnjb3DyQoDQvpDfaUYUVFHgA1ZeJqrcIVz4cw80hUVVMLV0aP1ZFM
M7P32lFzG88PkkbCwIDpV0IhixxYXnuUPESTKm8SZih74rkOdp9KOCudUXfvfL4rvGGjUgdyULQW
kHLWkriofNmjriBoXGiXypx4GeSNjUPpPBwruBtAXauEjRfhLCMvUCiHwxDZDJBnOcT0bECtffhi
SqoYSVUnT7X/6WiohSUpNpkozrbA6IFhukZXeJVfc3YsVlK28aVNcGSbhZwBUgZbADT/GA+nFQvP
F6nKuPceYHSVqx/ojKryPDxNvhZlIcT8VbuYhvWHxPxz+wvlwXKmSuXIotL5BG7nYpK/xORkqogI
y3OD+48RfDie5HdaZBOXnN1zT5PN6yWF44LjFaEFaZdTcON6RmGKg7Hyz0Yqobf2AhCgF4KaE0ls
c0aW9ePtbDBX88MMCDYnC2I/u8HLrsEJDZk+fT8JsCnNJPfBf92Uecvk7mpnT7Ai5YNxbiQ8giBp
lypoKc1RwpN99c3rv/nS5c2qfN2+RvdIyq6jPBCpO4Rj2Lp5a0UAET1CjfMQ9ukzE6JvtUrTh8kq
LrRsOMDr+EqMBEAfQ+i5LXjixjXoR6SV3/wrcU6ZbRJxMLsJZDz6jGqQZvXXqccNKQS6NJDqg+6+
Y6YJM8g0SOwgcLpBXCmEJaK3Hy3qOjyiLPfvXaKzffg8Nwq8IK8Crk2KUX93h2Ld0XMU2u1ZtlGp
oUYDXN3LC4Bx8JTIR5EonYtUodXx6niaBkbFQW588RrgBQzAcROlaUKjL2yrwmey83ulVVrzLhKW
y0nmSZJyPLYOh8FVU9CzV75H35Rl/AAzg9aqNbeZs1gHDqsCK6tI9rOuAtZ7P7RWh+vGfIY+s4Oj
YDsRDj+pp/mRhVJCamYdby5hOKUfRFE3yZwanLFAGpl+V4oCJuxdhD33JdJghUm4YudkLGEk8pyD
E2uZYk4qi5VIyglDjy6v/w8E+yOPzlxHdoJ7iuf3uT9Z/kxGwYJO7KHcRPkUVDKmlJGIc5vrVLmR
Kom2Zv1NTqdQnoYdacPt+diAEtgPcOR7NDHfnBAjZeIv+GANWeW7tjqZAfEFfbb78Nh/5K2UDZKS
tTS2fWvVh8zOjnIz/W8vT4qwIw32iwo+avy/Qbhv8fpdKbfocvgGuwtHUUYKF0NRzXH5XiavNEvj
6ZDo8v3u028DJBeDSW3P8PvYBNU8jZClX0fvxqg19iR4avjuLMt6TftH8EpUGVH0SMf4/gXj4akH
BkMTu+o4cNXQ48iuoE6mW/JeBTNNs3oKerw43WitDBt4ZDEOFsw0p/XQxODhbWe3/8ZyqywMlU+a
/0LudibcbFxTyCxA8pkNrfn4MqX/qSqNv80mJi7ndolMJJ2KcTf32YHicpExgDYrZlHiIxixurhf
f4U7OwHNX8zTukAcgJNgpvaCsmhADJDdDZTBMkkM9Zys3Y7+hlXs4gv1FgkXgcassU7hCgiY5hm8
19P+6648jUpYNc0xj035cv+lB9dTZs1bLZiesMnNfhjsC66e3Y4ro2PwQoKbkPj1CHfLvn/zP6wo
HTlWD95VJwkY+nUf6TubdPqTmoyAXhAw9WjCeHCoITRhniahwpi8zy65ntvqw/4ZwQITz7e5s7u8
+gNE4L6IHfxKfxLYVJJKqnFgnbwBd9UOrifh3OizE4WMG/l4ufqQZg6SOrY+gTtjqdznltOetw98
kIEAUOfUSWFetRGm9QQIAJtr6rC/VE9yW4wLXThXAFNLpCoQdrCL2SbCWCypwAPyCGFEHBKONH3v
4h8AMLcrwbtsqUr0+phfCa+UKEeGp7IAON1lteOTy3I1vluen7/wIQI4Yu/xneAmF1dwPA97j01a
CAmkPboNs7O1WZH4wbq3Wl7EOz62x5kQg4kZR4T4Ssy/ePuLsFn1ss01VNwdEAstgPf/gTOedhmB
7izIrz77A9rNL0HsmBQL4lzfogRIZAw6J0RZ8cuiZceNZIsUpmAHZJ87t+SH+s0UYW4aoe4dlAW1
f6hvzcnU5+xK5dhcqUCfGA9myDA4UbwU/GClsXiUZLSX2hwgthIiG4RDY9SXUIrGoXSGWRIa7raU
aKqw5RB4vOcKsksgmKKDA+QjOWJI7w131ySWhjPSi36SCY1vp7+rGWVKtC+XDR/yykF5XISbsAJV
atbJD1U0bVAxUPt9UV/Rckw52ozdOcSdZ1KpM4XPgwwGPSRI+acxG5ToWY0T4x92CUXnA+0DwqmC
HCa5Ieo2VUx4b6Sd3eoan0hZuLaFgXwDLWgyTqnS4c52Soen1zecrQhZ5Qfiw1MQ7c3wuZ8mucre
9xIN3hkxF4s/gQbldn5Sz7P0/rElUZQn0fuPRxfb7aIrRwp17MlXJnBJfk6Lol03O6YiYpxeyVJ+
Ze35XX5Psr9TYWlj4XuFfevmlWzkVKap9EH8BFyPennDrQOzDAL6f4B6KdgANHNnHwA2qE647eZJ
yl7CYkThHAnbEDrc4h+8a5lmM9N9zZLR7vBaqOA9DBbZ1G0eAjDdYbrmHBy9sywmtWeTDw5kyZa1
jcc9PYo1VZpwUVSs94AOeOWTwkplrVdHjv/ynIF+ViWlZ+RyJhGOOU1/Y4W5w2aOFBAbRNRop+ye
AnUkTNPzHKiijWX45qYbkgN2zY+KvsE4IJd5+bCJrykUrtcTSEMIe4Jwm8zlHKtLddSXJgGBBghr
O2XzSgn7xWw0pGDx2Es4CjTby1xV6P2aq7WAhKErRzciQ1P9iLw2vM4f6MAv1qtYgVYEEIoBiEmA
rsbnhvz5ngUr284EtALJVG4bUrZDfeOMv+JBPBgMhHyGUFQwFS9GoDWpfLTRRq33ZivKYJvmra5x
oycsJmxWHOY5uc7ZYk23FiQUvMBCFKYaXaR4oaGZG7T/PY4gPazUcE2+A/hpOrzJfyIlcsAcIGck
nqxZS/sc/WwIhhKNcS0zTXtQ8vAbXy1kzhyiPzxa2+E3d4aFCndSXiPtrMcVWMaWloPpON5J5LH3
y1Jd56hvwzcNMy/Xi+bFqwowNmk+ygNKv3fL8pLC62HkyOPmhowS3RegVOV1F3TmTeUBMp22i8vC
HAI0lVX5rrUq0S+ojOe538ibowosPXZYmGIIyqBby3911GsbtnDx7LRhhNAEvK0xW8JmeFxt5rR7
/CghIDOlr80AGvhzZwrGHaFc1gAaxbT9LPImGxGvxXH93gMbFrQbKUbkEKZKxNImQZstJRVvhHVc
Za1dHRvESRzKPOCbrknnL4rFHP+WMLAlPLK7L6ndWyQgI2WbwIQWGkxs4Rg7yby0+si4RdadMFjM
Oenmp/RGc9ydOnnjthudquEhps3wq+r2ONf7fi7ZHBIMSP2+zYt40YvQNc/UusBosovMm5e6DiWQ
wUXFlCC64tT4tj+9WpMe5xMnmbgzyeEOK2fzTruIz0c09Oof5V/oNv6/DQcLX5AkcpPNhcWuTV0G
rcGiJQzUm9r5gjGViX24L3Ea2LjPYlqhVpQPTzjXeTFB8aeluXlrxJHNIC0rvdqX0ZMkb1dL7cgj
eVuzka5Vvn9QqgX5GWCdKS/ljmyDdXGOFr1TgpSFdv8rpFmYhE3OizjFLMwjYy5GpHnWWOz01TLh
yYRXhCLE8IypFiAKz4J+zIzBh7huSFaaXDPsLp/PuTPKMwvKba7OZpmXS8hzHD4Me7hv8uoiYqVa
be2RG1cWz3+XiSyEx6HGi2TLYiVBC9PlgZR1Anw7RuoyghbetGSU7IwLjWz82VNks3IiYBw7C2cg
mx9doj+8lUmZNGEn7Cx/ZeCTZD5UfCNQ2PZee0gb4xWrHjgKejgNPwGsXIoyRB8fVpw7ufNxgSJ9
NuSVKSjwwtXG1mEaoRtJrjVHNBkLO3a+jkkL6apFDG2Zb442qOskgB3C+LdanbHmc+ozY0LJseZL
88L2zu8RRK+11r+85yGkOGOIPCjt017/nZXFgJIdmdeb4ompjgLUe5fLnCkTT+6PtMHlhWebItpd
Ot8P/eL7Vsy0rnE65fosE1knxSIhPcTEII8KF3O1aWUjDvd7h68F5nZ+AHbJBFFOM4ceDbGfjuMS
+8ZQK7Mr3dLX2fUfb/VyEcbhIZ14/86C7fMSH4btsDj2lc1xBqKlSy9PhH8id7tPNarZQaSfYFXd
/cx/tIJUdsXGGcV5ELP4leto+jWQx8WX4l5hMCdJhxPocn6HXkQocnus4pEgDJQxR0Ada1BYKjY4
ZbAc+DsozoZGwcO0YzywlhNXe+X61eb1t6Q9FGRjfi7a/jfVcV+7AIRW0At0MVoZvZeEfgcDZ9Y/
zC4vOZSc+kgCEZ7OBdAJyUwsF0SDzQxRcSBzaVL7fy1PyNkEGUVfwBOk7Tgx0XeqV+tnkA+5QTIT
g8Zr/Ob32HN4CZ/HoHeP6lOHm3iOru4gnPxSWjZ6u9NDUs2UDrrjriKBte/yHoHo+GjNcXVNIGRA
jq00utwQ2M3LKqFBtwpnubUEJTvFbsRN4bKwtRTClspPOUUpmBjM/FmL/r6uvyz+Lhn+s16N194R
EDTz2qv+eN2L5aNLCBbc0SbyEPm6GyiobMzaqd6dLiaq/GLwj9J5iH2KQA9mVvtx4XSi+t8VZBdR
J9RjupjSkfmAKIYj6KM6qHsDW0alVuKmbKpJJ08PM2OiDj0QqZMyALs00YCdLuUJaWORtPLgdaqX
/ydCf2bvRLQ0zqGmEPuNTz7gLBIPI9sZGfn0VivTIgkvu7iOPG/H7nzF6rJLym7F6+EDnK+/FfvI
sAde9l/Eh2QZNMX1/XPn8w8ySpZg8aiSQlaJJwSU24L4J+7pB0G6HwzK9hULYJGOQ8S6Pko344VW
0NRBjhTpjAA1alpIutQqKQtItCea6Em1okKfrtVaU8az9YpD5LrJe0IJGAKBjcLV6OtC9dgqoK2X
Lw32uI6DpYcfQEGX70pOMgFKzUa54hUMmijSU5ekv4Hj+phbliK8MYMQ9gUszH9MKri2ZmwiHGuh
W7Ege2xXDcle3gIeos+zrIGVO0OwVuCkCu9trmKn2URXiiRRSsNL/XkDQfU6jG5ti9lbVD/GxyEA
KKc/a6yS/rWgrn3bo1LmlbDIhpQ6QOPiviyhct1BWgqRgUi4m11PxFap9lfBsW97S2x0DjrdoBKi
FJd+g08QDgqeX89dyG86e3t2CTSDvv3xeK5GmEKbi8OYgIec+TYg/5c4JQR3Aht/8GoT9ILHUGJh
iy/N6qnu+Bf/Z9iOFo/7gAcBKXz/dRCgXblM4xao+TqEdJED3zVY3R5JyeQ8FvMLFUtQfOamBoMU
/1SESI5EZ4im6KqvUwHrV9Q5gAGKBkJvn4Sx+Bb4L8php1/pTRZWN/twy4dFBqIvJDiI898gikqH
LkC541dZuFrq2ZVYtspJCVeXeQHmZlIvOyZL5Z/F90ISXb5xNPJ1omZJUJ49ED68bRftqOzXkqWW
D0+2GZp5TzhM62dE80lRxZSCsKgSMAJuGiiIo7bcSbe8O5ZfUuD/Ri79rwe6zzTkGS7zYqJJsPB2
GdroS7dYMTbTDq/I8uFW3XtqIH9KTltRq0NOMBpUFs71efXwRchAWJ7lCUZVDBEhwg5LS33Gp2zl
Ng8miwgbQEXX/zbxZmnbyBPnkq1SW8neaxh3XD+6drTsPF3CKC6eZafk4V/76Q2cdiID21A3IIBc
ycU35xvG9cioG2rzbJPL93O8QEUDkep1qVC7L5hgGl67XwDv+6kNCoAN9Km2HhpP1SmdABCQtEyr
Ep6xlwP2XsEUcK1t7yyNWN8TsLOrZQcTMIiFr5EFge8nQ33k1RNOBoivBmRIS2FD/5cMnuGJSgPm
fRsVmhco+OTDaZDJ90gvx1AqarpvjrCc4bQpPG08zme8ChXVzN+d4hODp9J8e2ZmTzP5mmzXn6r6
+Lqh3arzurTtBGfhPyOHcNMPCcwO8WtLio+gb51WpmbfNkzCzK9OIMMmzXoDNBm4CI5aUp3/i+yj
d4RH0BIsYMQASCUmrzo+sQsbIIWIRPy1XH4VQNViZ7XnjngsTQvnTVvHKV1d/N/VyQHdF/5F9iAm
5EdZW9mho6QiQGxoo5TR4yiL3P1bpOmSmSB5K0IXCJCxYhaWFIprlBsnJyTeHLmPXC8xKZSX8KfR
2PAKo/DKRnDolJYyEnLd2JGn1hvZWdGa22OqvPWCZXUQJ0QGazOvXxY+HYS9ja5FlndoalpJw8ib
dgqw882tgJCodC/sHnNUaEqAR5B8mX63wiC0wyGFq3FqTxkT6o6Ug/0SNkvXvBupM4c5J9cZg/SD
PapkKPs2BjR+4haLrqWUj/WIeNG7LSYaSY1gdUbIAvS/8xnuR9A32xREJ1cHi89JWtov4gFjI7/R
4PGZMR1hu3m20zzWQYbrYueZ44WyCAiqQa/B4qPFlLkHcJArHx3Fm6kj5iSF5fnCBnGM3/8J55PU
5jTB8vPOoidMP2OoGJSCjuHzIGB0hAAC9+FmHImZz+1SNY3e7MIrxK36r1CtH4A20kdJGom4RXHP
N9Cs4ck23iBD6fCzm8dhlLLKIor872WZRQs3rIbk/sYdLOJjienVjD/C0djovtBcfjRpEXXCes7z
GAM5EAWVpo+uXAACodimLQ1vVTfSR5gszpR05ml7kHFEJgS23wDkwwzMUIB/H+aiRx5tquKf+CSr
dMrWdhIBtQdLrLMhZwc03flR2MS3yRFqWcWB7CVFuUdtVgJ9W2Om+MoC0IhATXoDVj3zSrg7xk/G
dVV+KWY8uIZqfWRk4+4rwxOLRojUT2XghqwdY/yCGMcYUsXwTCUEnciO866xHlvfdNaof3M+QN59
ZQ0Et0rRsYKSk7Y6JGen92+2/qeOm3ga+P6D2/UaSZhLnuSCSbwBlw/+UlVQWOfQWU5Dgytfii4a
aC5z43uiluMMvc23ApnbWaM+eiptrzqOl3+1es4Dt8aqiq33mQgtcD9dfwl5Myd4m7HP+QB+BDKs
POCigRqcqxrB1RZwI3o48cOH04ax1ibAqGEEAJm4Rnp2N20OgL1Y7EhGInBzepSVhn+unPm3XnJ5
/EB88b2fKKCGYD0ciWLhOV7bx+qh8ktFGptbQWKRYuWQhQdz9WAUmy21lvR2XrE9+s+PxaVdb2pX
F5+JzvuQ7Qz+w4J2Id1h0iabAF930n2ze53BVnDzc9c71VEHWY5J7fdoQL+l5U5gfv9pLsyYdiQs
yJ9JHO1Go8KPQ66r6INDr5ITETSOwPOn3Tpg1rDjffbDEGuOwEm4BboPkDoUGjSIFPq9eLpKmk0i
6rxDWC26Cqww4OTuJzwYN5OSo++B9Hh9j37Yatbg+zfr3AyEIRUdT1Ewvn+tgCiOIYOYsUP4KVyk
bmqYiTwgbV0JQOZwNpR302QbSuSNacY5gCdDbbtfRVLcemfcIwhvduIx9TkSOk8c3qlnp7GN7Qtw
5eypYg5EXcYo4CDkGCnhndjWJWU8nPqw7sSmKcDSsz/sLu17KhQNBkToJ2+X/hBg0tKlp4C/wjrd
vMf0nK/w3idOBSE4QsqW90hkHqMSIaRFRNzjAGOZw1sWs8k8RMF4Qdy+i7p+xvE0mP+81kF+8TQs
l+I7UKAgTrQoT+lZq8HeJCIGnBPdVgaOb4YDCjD2nyA3lwrPv/lrZSBazdWgaYGM3TGBYYMVSOzp
l0+ReepHmLwTTNmd2J0F7g7bogQ8/gu0yf8rK/HH9tXJafAJIzRLr8JrQm5P6ahuab1/eHMtAAE5
YyUYvdWR1coBSNOArpcth1xozVKg8H1cNNUPg8AdH1gPYtCt9OywKLyWwR2yeKaq/0QJhSj/EX5n
FWwBS0lQh4Ib2NQhY0xocxPaE37oO5dMNvdfPwPOItuvqxIwhIJKCUrTtraKGYfkYNpjScUkgkLf
wrd6Z2RYPYixvbbiY7/5bBJEr19LXQmOV6e8k3l1t3mg9bWpQAiXRCup9ICaRoLEt1gBwJATUCN7
k9SveQTIV0M5HKd5XajWryoGCIOECQCogUycRUU0wJMEyHoUQDNYsqNRqboaRTkPdaOnhjrVrjIZ
UDkrWub7xppYLbTmQBn9zI6mkaFj5DcgIYg2gMyVUsgPYyGO4wMr1diG4YuoXpRjGpLBBEqhH+Kl
FejGELK8ay4jcnxs7xBXj1wTUF5uIoGGq4hV5ct+oLM6JkscNptN47IGdSAGuOz9qmWKOiakOyn7
Gm7Oap5GmiGDNhPZrs070Lq8X0ybl4tBpF7scfTzk0vY8OaVj27jWJrhr5dHA1fbfAYKF39OFHx8
CDIjZwjdsaeT2AG88FzDngHS9OA12ycbx6W8qQvqbfOTuTxsfnMNhAjeWlhk25l/Znr5x0YCluOE
jc/crA8xBDACp55EuwK9KA9w3EBdPtWx8oEQvxnWhO4ZS9Siz8iZ9JIg5tEbOjTZE2s6jo3t2Rpg
HJtVB+qg8dCD6kK3CcI03EC19QwasdhdmQUY1EiLvtEdf+G3/otWHU5xlDfdJ1RgWvjdapcWO3+1
qUxh9Xcw/eK+xcFKT7JMw6rrzs5PgQ6EJzV0s12VrgyM8axMexnRttZRGIM3Yv6h1EQQHoIv2oNP
3OGcGUA7kg7CkuhVj2OFZWeYp2q82PHzw/PebBu72IKZ+NRr+hib41kKO72JfTX3kV9rmBr319EC
PhKAhYG4UVutiz3Pddwvbkkvg9MjIplIrd5uIYq0K0mum9qvf48nokbQUHPv0BcFPesBm8RfskUJ
DJ9wRgvhFGmDEXLSn5ZE/AT8mmr+r5U9kWUm9G2wQK35dejqTdkjCPVixP8gXiEGt5I2k33gBIZ8
VKCQspsDbpLj55nvT5sXLdY99gWxDxPO201V5JIgdcfH8XKcf2uzr8hPqm8n2w4QNDNTZV/T708E
k9aIdiuIcrO9k9QIATO8wBs1QL1XF7jZdcj4lPfZ7V0E8tlujc3at/JorMPOSOmbRkG3hLVZAIvT
ygT6uTrznUO2CNLZzZkVIMWW1LIiovQwlIKyaSj2zTTQLURiB1LuY1Wi1J8rUeK3Rs9kneF4aouQ
ujASRUEOg91FlfZeyJuUi13naQ6TCFwG6Y2eiUKfFPlnXLEDFU4EFhn5qJA/4BCqxQ0TdEj1Pwwx
OI3s0uGlZLb7r3rFNy4dseayjfFas6R+NpDTAGWnXISZQp7PMOjHXv24X+kWOsU5FWDA/HSxXMwa
EvBizxilBSkLVb2jrfxjw8QhRx6qPc4nxmPIj65RMsGc0eX9XAi+f1bv7A6V39ft1Xm3aXXbowkE
e1jhUF60X59HI+wIUZfmaJic1pkLAtYHC7V4AkCMLguLtxMU9zs7IlBZ7lFWwevNc6IuDkPeyuje
cqNcfcrAZoNJKFSwt9ilhF5Jp1HlCjbwuD8T8jn6XivmKp3hKRlfSUy8cNWpvVwj8BTnqsRFrjDH
zj/pfy+o/beR2blzEZE42DK8jpHyCEuI1SjWL4p/VPT9QcQhGlRPO+BShQ2tvZ6dIip2INI0at5c
mXJ+oqcfV1wN2L3izYBv/nlLsRHiH9g2has/HERGYNjJf+Vt6l5M0tUbmhodmcHdkXAOs4V9wFjT
mdpcmoNw0dMbM3U60o4fDp1MmvC2IeNC9evUYkYM5qwKcpGjlx3nCVYxyRE6P6ude1WfIjCb+LHu
/HgbKbkdPZ98JryM7+8zrdpOAoQWu/wuRno+AvRano412tPQ/6ujdFXquh9TpCvD3ABcbE/Ft3HZ
K8IyNAXqFsJC9hcdSSVzzTEuVDunAGMhBQo9YtSUsffO5R+bzruPrvqa57l7Fbb5OVAnMf8uLz2U
2ZkcqYnsCLAu2fap7wlcNfVtNPTDlJpk5AIuzLFwbQRKE2L4VZbeRK03EuiuU/8rr7a+yzUwWDRs
2YGTi9nZrW2fqfuRrLnfaksLCHSvNWyLJTT9Awy+MPfh9Vjyni+7VnNw4Vr3t5pRr6+L+NQd1zB1
Rm2Km3c/uuok3Go9inyLWUCTOHXtDHnrAFWuFpK1WoI2WVLKmy+uxNUkMBxKGd4suA0KaWGSN/K3
6Vi4fz1ZIlyfa1rVdAIm2lWsycbw7oNF6mppa9sLy3W+T+CbWfFBLWl8G40jTI56FnFAC1o5g1Fk
26nZh80ZraKCrMkovBkCplUn1UzvYvmTa6r8AMG4NoJlnPuPFscja+cL1Q+99d0IdPMy9wFfrw1d
NX2BqQc9zaLpKS5av7lUdD33zJ/emSihbxuKqAhs8La56EB+ogwMebRKYQyMkA59GphuHihdm6sF
zg50pDUdD2QLmE7pQFX/PvlmtPNCdDig8uQnFknirIBkr+W8HMcna8RSpFZWoylNBQ3HL9dbdknu
4FoU18vzrc0W5F56wfKxNVGpASkdd3gIFEKKjA/7LY23Eg1A7eHxo/mhJSuNjA2UyKusJ170zoWO
Z2XWtIPbr5gI1m7eOWKlvKE7f8z/d64ElfbI21w13bS4renU8oKaiNRTcYrFe5M7nOnihZx0Xu7W
hZyLviDIZjiyCdWEfKn0/a8ROP9foYJ7ycjcRjlInRdthjiuUg8oGT9J/CRYfblciPAuZRjd/gWb
LI/0L2dj35S5c6arthc4WVIH1GTRzQyTs5dW/x/3xQ1pFQljwjoTSbSnKK3rY4X5TmFf1a/JgF2v
F+CweUjyNNzEPQaKgx2XK8ppjEw1ZXt5/zvrYNQKcSmU2AHMMDH3RS+XJ45RpS+PDmsBdjQdNif+
oNIiRgb3nyzyccPMdKZl3KY398ovbkSzew84fk/H8H55LIiEK2g2hH4TlKq5GDpz6ioMFtbuJ4vL
ucevXp6lWTXGODSDX1LKNhFHRmyAhcw1c0PZeGA8ZlHAJnQ1H7GSV5qb2P9R+zmxnPpA1te4yq5X
Ri7ltSHncPbCr3sfVY3sj9fl3U4dNYDyHsyrLqC+9e4oyZaBAuHHRlg7Dbywu6xoWkIfHN22v1HR
Wn36SnPp+wyn4JnFF53IZw/T56NsvBEdubc7RBC+KOtHZaOejvuHNvSnUi/yp3E3wYtW3k9QZwUg
wMy+UTmLKuL5+/iqA7DVyYormV/eqvvH8ip7ZeAhP4pjDnBHGgnNE6EOHW7r3Qn3G3GDUFgPAOh5
mpLnwK0ujnSRxdg6pI6SFYv/6WAE/Fiyy4hRwoCxsUrUcgGgagHTJPrwaCb5S+GCC7Ju5enccB3I
9Rh6kweTeCZSWSbAoRlhEdtIpebEWy8usC2U73C9LbtbLxzpUZ1wP5Ep5jgyYvcb93WU8ICjyY2f
ALvv34G0woXmWQPhdJQ7Herf+Lra1y/dJ0TsbbKNFRgKZJTqTI/V3U0AFQ2MccnLKOalBILmAXit
nZNfrCGlrTTgfOKXm/HZBLVzqgeDxbkckxCncF/RidfIHUxQ4pZpac+Wo1NO0IPuhC9bk/Tgm07W
jxnCywyM3zptQTX2WuABjUcqDSTGB2acJMU3sMPiTUOksgLAZliK6Hik2pEQVUvEaixp6zqIm6NR
D26t9zlErzd1suVM1fgF47IMbTuWQPOF3mvF/VtesGOL+8maJIEIF+jMu0yy1zz84wlrGcMskLy+
wsdUU9tToEWSYQrSawOL48j0ay8Ou/g+JasHa/tcjL28aA8k3dawjmAisXVtAPRE0X2W09iytgsq
gMLemKIM7afxZJGVu3N/w2tGdA4zXqWxeUFd8rCWuH9Q2N27EGc1dYc4wdtfe3n+NkF8/2oRAY/i
VuZry8psLqrGgDjN1oV/cptNFWMwUApARIfYmGl77vu9Y8Gl01vJ7LLdv2kBEOExUoka2IccS1BD
eS6/8UC14ZK4sD7zibj53YLq3nnYW1P8xomh1p2CsGQKGZq+szoEAwF9klBKF19aNsTHT8NBMbhf
szBYOxWQEps/0nZj/Ti5v/9M7VwmUOWDj4odSe5si4T+Z5ByjHFoVfUewRDz1FcVWCKZ3uBEQukQ
MjxFW99FUoSt6MW5RtvsSmiEPaQn3vFUkDT6EW+HClD5c92b7AjMK2LACcRGTEwXuxgpu4sRf6R9
7MZNWNl7rCexQlb2BwcFyf+MitG2mCLsjPuhafi1pEk58ojTu5ahcFV13XPhh/QRv6P/sOOtjiDS
PxDeQk9Q2uQloLAWBf6Rmyu3DOa4fG+MJHm5Bvv13PhTJFC5cSN7hAMf1C9xsy6GGkXMQEovYNk2
RGHBcHEmOJVFt+gK/kxjysh+vpsYp0GQa3btGRH6KmeVVDwefDpHAOEMkGC//NTZzgk/0K/b1eWj
sLjfTIJDkHIHQXXfM9e6rzUfBYYRzcC1tNq9cGx4P9RRrQGbACNzY7OUTtKhRrcRA4fB9QUVy/UW
ZjkSXWl8wmxtuCLD9LRDvEdmhcJs112QVuW0hvzkC/po2M+fGgYpn0ZFx7pplRg3bDWnWVbEqX34
3XvY0I+c8iz09mRKettekr9E9SdxLRkNw+ME4uSdwZ76zOt1fiTKmQeLaHpJXXAvRYsHPGqtQ7bE
Pjm7Gws0xCdv7PZeSJ6ukg3wkC8K0A3F/CeHTeRsD8Bev+oAKvwItV/c96JtC8A+8YSVz/vFEGSg
VBTZzxW8TLiWY3IeW2TNPdkw9SyaP+3UeEiEYtUxd7tBPkUpEC1zoORiI0nw0x7F3NDcaKd1FtjW
KEocZeBUDPsIhXTIEMyk5epFpUs62d9cq0FSoPK2EAe1vr98MpC1Nv2O3ypTdMOW/wkTLVkP9oCE
9r3pq1G7c1D42SxTUqoOQI5n2Q9TV+WLC3PHXBoVspnCPvpp6ni2Dvl/SoZkarkcUxVDe7+7k9si
ZWQHsfKy9xTuVpw8ShIxZd+BqLINflPzXShTF2OqbgeTGqaQXvwCrArNguKHREZId6Ut6Qwbe1ce
UreWk50Ejjqmxgcx9j6Unb8aH0y4OY8CTktUqS0wRTDdfYuuU9WkfwK7t7bKoKTNhgBRAqTCe0PE
AXVUui6W+OS3HSIJ8yP1e8WvHLlusRDJIlBYQ2LVOtj++p3xDHeiW4G3kSQqMZC6orfrxTrqrbmK
CVa1LyMQhyG+dtbUbAJCszpWHpfGvwqsok1M0MVjGV8OAUG5UsCsgDHwhh6fRbgzrITOhc1guS2O
jPG+RyHXgL9b3CHhfPbm+q5jEjG9opie1zzJiwRh/KU+4ls/cc2e9D198FOc6Xi5gukcu9wjC8ef
iXmCcMYYhLjIcC/czTBwFhxbv9z//fJOoGYPFsjUTINMiVyIzLo46U/BJaj3ASMtwjYGwqne0TRv
9oVBFWGxPmqJQoyiffooMf36a6y191ejoFh7MJAB4+xX25pdkWdenz+q2YIf7PeibRPR50vTeASF
b1cpkS4Vx+dLuFUbRmXq9mtoYdw+r0teGEP6cs1IHkxL5+9Uq+E4FXl9Jswwog4SU5Sg+tEdWo4A
Vz+1YWZ7DftsdevvzEH8TMZB2VHZ/CKG4e+kkac4xanVh554dg4r/OFjTdKMkkOQKpvFWd1J4Izu
5/rxhH9Z2r0oxi+KVnyCMQU1SypYuctP+1n0d1Yual+pnv4eS9ieH/Oq235a/+xDETQsLq8WqGrv
jd6XOFQEtdHt3p9MMvbEb6BWgGY08I/zPzKnO42Lhi9wy6Km3EXNJ2IgK0Jx7ki8wrgkd0ZE6clP
bGcN/8fDr1MSqQFtazKfVdCchIgb0+/fNTv0bvL5ZGMC6+0nIVqNwl1tkx86cy9k8lLLM1xn7CQt
U2wprWKnz72HQ5MQbQyJ8uJzKJR6Ex82NVF+nANvdk69PthIO66+RCNjaOIRb7VYGMEIOlwcw+bK
RiJ/r1xKX7QB+5iB6TBXNyBh5l+CDFa5KieTneQERS8izSnaIMo/FgUtQ3cZ7xubyUym/Ceyzf5c
HRRs4QtueHyjPNElcTs8YEo+cl8GkD6kbcReentO59e0FXPJryoXbmXNyZ3C4fC3BWoGSFjhAynI
AK6ZvQCJRr4t9bACUYw01dQMW6BZfBKmAxNchxqtjtd7iZCey17YaEEiH/Ibeojmj0YJM5TkjQpS
OB7HOe+7ECj6s0mHSkOhva2aG8/XiAvr/xU+MDESFVYLGS/Z0lfZcw80KPROuie4U5wJ/2J1Ia09
V0u4LBd6FdQMqV+2n0HMGZcsuvVGFNBVrFIQCTV7UqqDMpzPHK6ADtTkANvv4OQQ1lkB5Z0XMkNA
kI9GxOKPwCFWpAlLogi7h6EHUL8M5tQfMTWA/waTHCt8Wsa30CtRu9jMLJ1Ax6VUMCghnvw+Z3Ge
V4GKz/4UqAlI7GWnQhshIJUINan9Aa/xOjS8RfKAVknwQqE6wpDHh49MRCaD61+YOsgEHXTOEV3u
ZrN3insMe4raX+cDLF7rfe1fp8sF47pC3xhqHv5EbaBEBh6xhP8jRXvMWjnUKXFolUWBVWX64b+B
YCmifDVo5bl1sUs877zBeBm8zwq04C6QMiwxR6NB+osh10gjqK8aT7yNrlH0Zf5Cfi/b/2fnQXL7
KT2/nxtbbuuo0vl8DPPN4+X2DAW75siC4miY4wgCa3thAkjxMzWh5v2cTDLwCHcCwojX9tomEoLm
fLINuuS2VshUgpi9vVdSHHjXlprIRxd8CSu8AQ7SsYh1DORZ/ZkV39J9bNg/aCc4jVN8LF4uryde
QJsJhE4rIW9s6NejZj6YhTC/IRd399/F2jYd6erIrmcqpnOdbaYOFEwBx0w/Tpo0QqTQC3G+QkBO
dYC/C+hKh73dNLP5U0phLRXQFXM/W+jfw+xopJ03v4bMnSpxrr3sRSEW2xuCE7VEsG/NcqaK/IOe
0ajrDfQEzR7mZ2n2cHzIwetH+2xF5BPaj9eQMRfUxKEai1/3Py0otVdYZqoOhwW9sSnqykfCJWJ6
Im6ZiNHUu8vUUlDiJztKe2L9AbhuNFPsArPBM20e95xVg2v2uMVsYgFoGHuyVQL8kV9n7577ziq5
PB0+5EDTorMZqHu4U1cZhbmtFJkS2DaJdSE0Zi+cKetpjWfsv2UgvCXBRsvwQjTdLN94L9waP39E
iZl5Htesd0wEui7UXfVRgNs2byXYeq1joQY5mH5u9sC9F1RfMfw3CQG6BQ5MUKpMpuhhyD2oV/1z
3nWaH9TNgJlb3U+JbYHKaSmaxU5OjzRxCDL9QxWPJKsZHda6zadhPRNRqqptoJqgqWRLFZs2J2hW
zYAOdjb3yR0ZXq0G6O54ZMh3d5UwdXxhocsotUziSVdqgoXi6dXGdbk85mfPIjP6dBv33pjm6WMT
hAgi1mIaNA21fPHW5Os0s5GqS82Sl80F/uXdZWR7UaVrXmkDekw1k8GX4a20omWQZaXHcyvTv9kq
FJEPLcz224g8C0qBMR/KoVUO5sBtQjzDWeO2rFVcnu7qLeaz7eb0nWEG8LzL4c+yFb2cX3n3TRjx
cHI8fwZ8LXycDD4D1HDnheBILLJNXHEMZbdxkNAJfCX8mP0W03Z1Sr9uCFL4ll4atm0klzMwpclA
r0IPtePC6hw1rvNIukzsGpnTXt73fHj7XS4WVzxiVvEErgKoFjQnWA32QGU1iSalwYksw0aLqeNr
dj2wC5Lxza2gp5ikU7IGtONFO4OrjVBGZdK6GYt5yLzk1ee7NM16G3ROJKrEyX+yImLEfYD1u/gF
NGWtSYwiUNCEBH6RwuKmgsPVTsbSN1MEujNDCMt83Vn5bdnS6/tWeI0KHgRD5aOwbMaVGTW7J+q+
hUFspEVxNXwhRY+OtWigq3JkkQR3vF1e7hluyEdK5M8opn78uaIJD+bJ/I4YG1SMujFpZufY46Jz
U92KXyR/034Zq/grgcLHn85xG+Y6dF3pRBNBrd4zcSupsfu9fj4Zweru0Wxx0dotfLdwO/4r6yyE
1Z+5osP6XwK3M244E9vnzZ2uWAWVoAtV0v0UQWQyvgeqR8pQ6XPyM15sE5DYJbrsDNX9+E/8zbKB
k/64Mx/Xw1RvngTTVUSUTvOxSWAclpOquWIOs7s0yr8P6GQtAgYeLFl2lSnPEE7KjfOu10/l8OaP
Cx1WUqOKJk1+jqIC7/lm1gNgZxrROIRMrEw9TaT4dxJK6q5aPIAlMRUHc7UFY2w4Du1l9XnobHZV
Sh1RVhlryVRmg2sueJp/j6f3PRlDw1D553tI9wYzULq8KjmX5NrqPlsAFRcVyJBvxqxzOZeJ63BL
/Y69uiHzqbz/YBjPz9JVZ25dEItacQKj3IC9BcN2APxHUCiYOsz05/8GBjpUuyM3WWKGmPe66o5x
g10czfmcHvnxhZgMvubptwx7EIyIykpr1WUMsH2ZmvcA/pwJKrZncuKcqcFTp4O9gox21Y/Y7jlE
BZyW67yrb0UGqJYCouvfYeHpfspq7yoO+OVw8V7ArA/lDhMYRUsGTuSksCEzsV4h2bA6kFRBD7bW
+0iP2C5n+KVxyO7B5EckusOt80Skzq13cxr6NComl99oxFBUchKXEmZEMirg417tH6DxnMZsw8+/
hEZvq31j3OQhjq3Ct9R+hhbv2o106uncTqkOrkIdUxJYaAv7luliNZg1eoXjPEPZkLd9U3X4XSCq
DCzacMx4+uiqS8PsiP65dzyXeXlhdHZRiOgNTQaEnMXXhRhuG5Y3sSIUuY5GZJe0TxrO9Y8ZdTf9
7efGxmNVfPDVABrPbTFReGrz+ux4bxgpZ8MbJx7q/mR+tykbZn0fbYYNepNVlY4Qh9JFhbq7vbx+
Xxc04HToplhZTx/x/2+VlGDNtcpNfMmCIswf00Cxaz8exscu7CoK7xFboNlabtsC3pTa3tz+l1wU
mRYWcNTocNNS3EugYG5mdT+Gs+OQe8MJw5C18l94jqOBffh9iWsXwkbt/RiOPjOVdI1jnUkv/wIO
CQZIgaETzx8PqcqWO6s3ipZe3u7wve34NteHcB5Ix6kDfRnqvuijn79q/AowOdZkpHpPlF5dCs1i
IO+cCt3WB0QhKN5Sg3732M7/kQcez3hITHHNR5Z2CmrkUn4TPzfjRPDwHKGuJEL94n7P1qLxTw83
mqcuOgB1CdF46rG8//ozIY1f1poN8SOrjp641aYTvnGXN3oF9coytd98N5uNM+oDWzujNcUI2ufs
x0hRNQ2towKemyB1K8oca9dECGJUVT30ByZDLbjlbxSNud+rt5u/4JRslnWcSK+xHgiTpwMNMgMS
n5ISgcSz2reJOWtR71qT9wwPbALjhqx9ODaZvQ9kIosVdngZfe5dy9Z4FEtXi8pt9Rae+Ai0TU3T
sb9neVXrXKINf5ETeDzGtj9CzrXaBVTGMeevZ/ACyW+4Aee7B5ioC0AF+fjH7AbTEVPTeon4myK1
LQsqsfXwMbkmiO1N0Kzjf80goYZ+hvRYH+u0o4GxWrpnEK5CYVQoFXrJelRbqstW02nZfy0uzSda
ktsXM/EB6ZKmkUbDHmMiFCR+3FTa6BC623BeTDjSkgmb7TjENaaww4UIdtIVk9LJIUbVvo8Pohw0
bKaVTOZE/LLvGt7SVX+Nx7rfaQVMSPlqXXJ1WyZGZU3WhKywRdNxQUXLNS+g71mVvMQqNs27hfm7
nvZnIUFkCDStGqR59noaXo/yCAQdADtRv+1MrIR0ERun3sQDipe7uAByeJhRYyPkXNqmFluARsSn
O6mNHWmMO7ueEMi88XuVcpsvshMuMfO6GdAVOkW3YMbNm9PVui6vT0AaloreUhmfSPe8o45j1rFW
BSHTqZXCNLM2cVY9funOSxA5uzlt3vxHn41KxXeuMVv+bF8MwzSpHEvuTlwKf0VCcZW1jukD4euq
mciPR/N3mJ/wKF3t3pXk5D78UEPD3roLGYnQn/MzxVuBJ95esd/F8jZBpoYYOQTwUbOpbrR6KBMo
CY/XtzRO28iM03RBYfibziXRd1QYHvcIi22y3u2otl5TnSqP3N2J63a++mjithA0YCjJezlnsBbd
0jS0fvc/3OB/Srf8qYl9nO+tt1ciJ43m3kZCJ8+soGTUiaICOhJL6wFkonerhMAI9rdcWPK38SgY
r8LFM7xT27H61+9zA8fP9Y7aB8ue3oUIV34CG26J+nnbuk7pvubv32KAI5mo6Ii5JaFxjswj8oZr
IAM81WKHwNArqYF4ULf9HWd9t2t/vz0hEo6F3HzuFAxA/sRoOc0ZUrLCIllQJuHWpjL//SiDRSGD
k5Om7YbbIHi9l+ME5cz/EAVecYAz2hOpaxx0yn7N+X+6CPe55eqBUpok0ym0DlDNitgjx/3PQ2g+
ZzvBe0dSEc0vJzb1USgfvE1u+LwoeL29hUqiTPmn99COR7WWh9RsvdoGHrHV6FIi8zAzm5w2LcED
3+x/MgfhPJ+NW+HZM8HcaKWWYh8tVpEJK5WHH2h0pBYJWcqlLyRXpE86cORWmroIl988G5pV4NwU
tEWOgeIxNFOMbOjIpZRtaAtwZsWJC5Griw0kh8KlKrYKgYCrSGgvLngyrCj3lWHtOzny7q8uo4Yy
2SHlkEqOvfjxaluY4hkqQq49tkG5t05nHW6kCbhpW+VgcQsPHTSQGXsGSV/qRXSKQg9tiCNRNWj1
QQH4oDB7XAqbeUzMpioJZtYyUqGon1hGalUqC+td7SQpBHFE/nXA/azfYO3ygOeuAFEvxnIghEA5
JgR4T6QANBpI4EQNa+IDmIub3pV8zn7UUpymt5iHsf49LkvvoNe6GyRuNp327oo/olCBWqf4FakS
HXaTZW7MXET0OFGe3TcStZKXZl0Tu92MiibT7ezSRXdYVqNT7NExnqqwvUF/fcs8DH71OViRX0sh
3KoWzw6Sb/xsPmg1nOnGqPAORtIQBmYg0wO/fkNEtNsyNbRomcPMHuIztbdIEu0RNWEuCXTxY8hc
QRPKa0OkHunp8oaFVYqFDaEgKUnCHh5gOA5ftPukwxzyS82Xu6MEYFV+uK6RPe0Bd88mwMQTiwkU
y9KfLr79oMtDnDOU7NcO/V9VqWkx3KESv1R8PUX5u4kQZEPyAFFxn7CfZylKXFiN5deR/oQN2Iot
skuIRQIhBHoBe+j2oMY4WtksHkI09Ta/G3pv38ougqyGKMm60e+GOs0L0ZauV7z02lHf864iVmWk
nEmw8HxPIqiQD5AReQpm094O0uXxpvbCesLWdkPECOojgroXD/9aJ5WK4jbJW91rrGa9QEbTnlna
wZ+BWB/tUBWgdvjGQddKxaE+hJ1rgSjBtyVcp8MDFGRQWf2EQbPM11x6mf8z9cC9QQKFBjrETcDj
Fv8/rVKRys+Pc7GSF/ccY5M0bIFVH+xZvxN42SZYLnzbBaUSEPIMQQMwkRcbLFaUGxBzgUJ2fjHq
ZJqkTdfBuwKYsowdhmUtnvELt432q5WR35TrnNbJy/yYjF+pCtnjrsegzXt+erO+j2Jib7qVmodU
A6CmjIw914/ilylowGIBqHTKUGdHLf0yQRVQjxAyz4HhlpX44PW7RngtIrSA+0RgAJrdq0jN0Zk0
SzSjeyVDNSc1qAKSDethyG1Ya1+uonQFcGLWiEfXYS/d1VNxMUm3QJmrg2kocQcdvmZ2EP83joqK
LnGFFJmIS29Q2EDuVa5GIoUGgZbD08yLcoP6WzNCZN9XdtLFcqhSSS38q+GFrCJfGZAQjnJNfkDE
x+CT+hNPR/0AKJg9xlxBNyvn1jABAb0bXvNyEtebe8Xez3N+5bWtGFX02NaTTyDKbkD5e5D3OPjs
A9zygIPLPpd2DCmv/0dXfvA0p0HoAPnH6N3LdPURU/U8OUMzsz2xFikUITKKq2iuLK5Zg/8y4Y9h
8RoylIeNwzQY1UsipNbHBPYPS0bQ62ctc6bjRquH+FV2lnK314mRs59FojS5FvZlgi4HgS1280tV
SkpcwP4UKqkuOsnBL9XyR1TS17NQeyIdepK5cRotAt3jJuYggEEL27L9qvapbxF8DCea+17SIzhF
Q+qpZEfJCgsp6i76E/Rd/3vz5YMpZsaqfU5l13M4al26uw48Y4p66g8Nyjt4KZP/UTBhd3iN2rZS
PgsU7iWRwu9DYKleu69Ips+UjyWEgEkMJake8KVwNzVoZOyT7PZp2hGTLT7uiVmtbQQSfdYrHI1T
MB2sYDnC2CWXywS6GNnzax1KLYATiTZjfISjwv8Ct32S+S+/q7HCz4j3BR/gMKPLgH1qTRgkRNV5
MEnFItqs74f0fz+LESh/d19lZIe5szkny0VJZO1NWn43qSblQFKiHMBIdNQJ6mcm1IkG6tS/Wx7O
Lp7u4ij9nVWvhEzRd0mFXvuHqJvbrllga5obLdCBVL+Pddb/eAuTKmAdyr09Q9QuslfYi/x5a2O0
6pGcCuKWsPUHg4ALJ4eeHF7hWxKH9NcRwzbT3Yp+xbe3jodxIbmzk1HgrqzI6V86YDKbf8ocNszZ
kjmF1HGSnrzceX9Qh1y8qUWKGjZhsHOLaPRYmGDTpW5kg90jtDSEpgR/mxtoMFuk7MIn+JqjnPjp
ZjQ2bNb83+IT8wx91UG7BMJ1jrUFTgGkdkRoKsB0jBEO0UK2Ig0guEUf5i9PzGTShVMlrTR3znqe
LqQJwu9DU6U/324SV5GNORAo51lLdcFvIGwynK4XdofTYb841keHR5cuKxC9tfCQSckHa0PoiYUl
U5tuvHjSFMLpH9o4nGpPpVd+tY4npKEdzvfdFYxZMO0dxLvdKusQF7Y3wndJTTVPaWoBtWHNlTT0
HOAogLdhoiRM12eEXuppMnB5Zp4V7tjqC5DCYBO4g6ydhoayau3D+kqtiKYaEHRQFy6hpobC/mtz
zcqwGjhqeT2lBSnvKe6z6M4f8nU98M3lcPPLajFMglYRwVtFCflhGp37cgr1i1qMx68R+OXuAiUZ
Tlgezb7usgZge4XuU0ALMl70FrW7MuTIlNsLQ1Md+sn/T4FrvIa+2HWQMvpS+jk1g6IBH4VZtULw
f2p6dv+hlCV9K576bEZrOsONoZlueNLtkY1iy9qxkRn2bsaMR3qmm8BqZiNJQt35Iq18FqwAA+UQ
5YROhFD0i3S9vq8qviEJY/D4vW3zbjHdx/SRXSlWFjjBUk43HD5g9B1dx+UeUk78Q3CrvPcNkpIR
4lREJBNvEp15wAW0WOvJ9q/QWSNHPRuK0TAsdqGK2Y8dyYJt1CdX4E0bSU7cWPGxfkuOkVQchK7q
m3LvpjawvQI0hjuLRHR8c7+NlyfyvAmRG4dUHf+nR/vKxjtzXy2iI9zdj1MWKKf2Vs/WJ6nK0TQN
e+7qDX57GtgGwSODlXk9J8pfJ7zf4rFORar/Olbyr3lLYOaNMkPd8uqCz4Jgs6xXijIrmYhGDBY0
il8hyXas5fPqmM5M8Tvi9eRk/ZJRW9Vdq7uVNGGzJB9oxzcqFle23kLa/EOz9bh7Ee7qhBNJaWvU
c2GD79Aaf2MkJ4nMfa1aUFy/kZt5RDZ5pcFhC6BWQi1sO6FD9NHVzDowBRTPx1hqQgpv9ff0NT/M
irLmp0+kqTeTtJS6kxgGoNg24nr66p7zFn9w4F05O80hudCqpDp67Ov6tbQFOMQgXcLLJo/FPqT4
BoBuMhdMwoeWrh3TSxtzIbax4uC3bIawANR2XS7yF3C1NpdZCMUn/dOXqFfzu6NhKpCb1LKE4h4Y
tWkjMmUeb3wqbXs0Jh7MBb7HhjJO5HLwYLbIw4RaqeJ7I1CVCJuqcDhUbTKxwJerW7E6SQ4/rDKy
RgGocgWyESB+SX/7DOpr6a4OPs/4QdLuTaolh/h/5TsF31tMYADpPdsrDB6AnOlwlVMVFlz5pi5D
6E/RHqHkmSETxrQCPf49hsXt2TR3F7/uP2JLcl9bHIFQiXqBXwLCqfs4X3O1FOVqmTkKk6XgmBcJ
Inq2iDutKC620Vtn9iISvZtxedRtH76uhG9VGLZjXv4+X2xlkL7hAfjga774v9ELTk3X+4JRjKbT
ty5wLVm9LGNmHbm+DlY+hbTIKAbF1l8EshH239OqrYOqr+9F1TQ81jdPLTgzLsykl5Bt4hiVeuFD
SqSq6EV40sucK2LMCbH/aqvzK8rruiICO03ByrlWesY0+qpoCmZhMPtLjGWYJXGq54/ruuCYJfVe
d63sLN74kA0UscOOertJUKf0V4gjj0Y5bJ2r/b7dDsItRNlzC/KtvH32mbCUCSRqbrIbKfXFHHlf
TqCdvrqwdN7fPHGIA0i+hETfpiNZe6Zi3C8nvgJxJDpxT956Uc4k/p8KM6qohVmwndEzKuZ8fHZ6
e4+jfgbQ09D35wGK/dX395q4yZPHqwc2d8+Tn4srqUjMBF/lSCNb3FxCsHqVGvNh36MF3ubbYHr3
4p1WCXYyZ2eWPM9m/DFX7/NZRGj+n6FpXL3IFtTqgvtv4xj8ufeEzzkUjkneb+4guUa4q58ERL5Y
8GhDKr/pisA5RStBJTACeySJNLc+qXBEQNxAG9I7X7tt2/FM4mbK8iM2BFTTXOKuy1+lwde6fAwC
sWOFSwq/lGmXyylKPkqeGiZdaYaGHp9/IkNktUMnVQwWiPPy4ZAE2PdbbWWn8u5zyhhdGSKDpGRj
Kn6EdTz66ejk6TwI3EAQ1d+frSIuyuqWncgoE3UVltqOfafLWqRiAYSoavANj+KlCkiSeG8YjnQv
91loFhTNiReSUHOut1ePXET1DLkTNfL5ef8ORzbb3Wlhx6yn1tJ+HQP5L+/zNZxVYVVOQ/Oy9rXa
CxVcBEHMD2+wqhEkzdf1wSQWO4VpwdOCWxmX0aNHy/9PuKjTnK/8zuM+/KiWzPVyX4bPcPSA+Fzo
plcrys85Xx2FgdnfKOvEC8TwjFHxRczVkk3xPcSgW0D1RtWSEjG3oub6HPBr1gpn088vAA3Ls/Vx
I5V0FcB3PmwHTrF2DVibJkUMApimT00TjG23Nnf2BClYYwv1gX3JlCfCVf+ng8AcL/t3T5a6XDrq
7fFBav3zVJAolHISvcL75609jm7TGzYuTE3iB0FYa/y22nm+hY5uxBCFntl0Y6rmOuUpIt19Ey5z
mM+QL9zUWDjz54RIZlLNSSVSvFwtd5JCrf+gip3q8qMOL0TtfArQ5nnLR8qy+7a+h4YUaiFPHLjZ
bk1MCW8OyKL2xqJvx7h19XJxrcSPi5PDmgw371X8ezb97gLG1ah6BCvTd43vN7iwG0mAoTMjsDvW
5bqStV8rQsDKzLOabfB1oZLwQbuWTDdO6gAjei5GJ0XlZmiMOr6bzfl7ilVnjCVtRETVEEw6pq+P
qdXtrklm/l/zA4ZOTeHNojo9RLGcdoI5+mFXnmUGmlGgoy1AifB7V7xPHSeHvyNIkUav9KZn+BvP
90UI2MSYJNP/L87fyHsbbPyVthwF1Eed6t5ffyLYk/XwCkyJr0XXgeudBUOB4E2IL9Ly6bHwMGhD
Tdot735hIeHhQQfYS5ud2P18LvUQSrU44mvVQpR8/0d2jHrB36JIt0lXRDCBFySBD9k5lVgok9KF
unhtgl3wNKMmKVGoaPjh9yfkJamkdS1Lo1heUSJPt1HR0R4xiuMTWPtMcOnSIrOL9LVDcv1aYEPB
kLnpkIj/AqZ9MZxatUsQZ+tWNBGCOlUl/pWSFMvxZR74FmN7kZvOvYXHNPhGjIUg1f6e5kFFaIPG
NkBJZ5RajB8AEWPMqLdbgMAuYMWTIE5c8Iav2mFMorHYIWQ7+OLFIq/cdJSypfLaHLXRSDofnC0o
BFN8yCmaptqlT477JLiERWjUmXRo8tu961/R2Kf4Nbi+8bZ/KTSOxoAqDdyXlNoBjACFXdUbIf5A
MQJJjYACG2nXNPXz4GYJPCmn3fvCMW9Z/ozVI3++unOfHa08cMn4aOBN6K8J+VolUMUIM7wopeW4
mMutf7Q/mDAm+p3LEUFtQDaA1CISm2dfZa76lRO82EsZXvYsmVL5RtxeC4/CJ0WXs768QAgmBgsr
iGimei0eYd1OvGI9sRbXuVUhAvHuEbsxfBrdx+BcDb/4+GIpU/TOtg+hIfTNTJT8bOtq/MS8WeEb
eSD3K+cQa98n8myCjLGEzxbTqWC/FI00NYYGcni7Zrnvzm+SokS74GnwM2TxBk7F7wXJ/J0hpvU/
Z66Ba3nCax5ISEl1RPr2exZQcDMb3X//J32F4ryQ6CVR29cKqn9Xdn6QCPtnew2Bp0ICHg3GjgGh
r5+w9Sd6mMj59V99Mnbe4LFKEsqeyvO0jiGnMXfaGqTK1sFOo8cidA3Q08/begeMAMC903Ulq2fS
k5tc+DiH9+eQur+W1wC7l9Yfk8X17AF04hsptSNAmqTrWJUi4wBuGLAxGJxSfm0w4CRlrOuWBEnk
WfpC6VGwdlJv9iqcRENG8KttBXveaeaE1m4xVkW0mDoXxZ6x1HzNZjQHsx77n6CerkslMz+y7QyH
HPphnvLW4n5Wu6o0osMjEqgv3Gt4SQvZrdPku90c0a13whg+11ZcvA+GWkTDxU9cYgYpQKUPUg+A
GdaOs08ORGMF4sUrMS+3YbK/I8FqQHDrod10fw5nX53GsfaqTEMzm4PYgO5rG3n6dWHSOyyVI+rP
wMxXwk7yfSMHkuvthX20fPY1xcGQJpw2A+U2eEaQHwyZ1GadHnzffRUKDYCeIU366yx3vdENKu7B
pqf2rmfKuq3Voal9VxR0f38IemOrApZPFJazuUSKWrlubt/kLioBk+4KJ9Ya7Bam4fT/koT0kqgi
8YIj9K0C16Y8te9pblaHexXj2ygkdo0QHDUrxt+5ieMDv//UGj48+2G6TNyzHzzxwya/U3fsnuhx
tXKmVza1/gbxhLzmypcxotP/wK/ahgcgNvm4BcPV1iw6YvVJEfuynTbdAmpO7uhCkCKTPcWArzJ4
OB2lOTOKJt07rnjKRlIYjmSdNSLV6iPMGQl5RrYPCTRD/JYRmN+5NYJBSrEYpzxbd9C/gmE0YeGw
nHQ6xspISW8fkA/X3gyPckwzjLV+mmoJ9b/AsMvJDw/9/4jY1gyiUHKpC3xm1JlOUPfBCbfuu6D+
Mtn4t6q9cvmwoR7BxvcmVSjy7ECT3YzRPeJbGvbKlfkJUocAb6LNwAejUDq22vFqOmCVu6O7VVz3
/PcueR+5tQVc0qwoBuJCKreUMwdDyKX3HcVRfE2mHvhJRWD6prkuDGCpJgdzC/dkqsCTVqEBK8Mf
QnVM5jXfJEvRdic9nQ4J37h6X4wVmRd6VUNSrXU9xDdjkac0Vc/VeebW8occz49QAN20r9VZ3geM
9emShUVajweyLm/+78/4vyXMztEszbMnO8GsTcyucKXZ0omYmD3T+3L6EH+jSMQxCi+p9ezpJfx3
j+glrv0e41MQfUdpVEz79cO1qJ6DqbHvHW8E8OxF/kL/+EV0S1YlIn3vdTAfYWE20qp+z3bxEC0/
jTGSes37C8P5wbnj2F6ilOaV6E6GB13ToN/yXK1VlQJxOFictEqhj4bSFW1t/G+7r8vjiTr2kyCH
3wMYluiMGHq8qCdx/PQL6BxiTPDZwnqennw4qjL1sD1QB440YdsOfbfK4dq/uZvtgsM5c5rfJRu3
BvcBHtOSlEOBqBGEujq7g/IkwLYBb52Ux8z3N6VFiSN4TijTsjr7XvvMRjrv/UWQ0J8SRLqRnZdl
lRLwFwz/QoN/5n9uzfFF0UzbzqrcW8vXnss48hrguhSqmeQBx/YbzXzZlFmVQBehIcw6lGHug4rX
F1YqxDkhqIqgm4QXXzfFruwpElqn/K7wPF3zBvsOghLSO20/nblWhOoo9ZN53aQWLgX873LZRvu9
tXkJjc8RpwJo668/C6oJnQ9xMLja5IbP2s3+cU+OMJ+IodRSTXjIi5p1gArrjOsacw19UQm9NGq7
OFzlWoGiUJZ9+VKUY4zHLlqktEu6OnYcjEVSVn+GTft07bUAs7lUXZ7qPxJ9cEG9YfABNvxLff/x
0noYJo1mOr54enlGaRYj6JwnV2Zg0cikQRyW64TWT6LuPfa0DlKCZ2haM9gHHHbN1nVjbwznWtoL
sPAgpgX5smYGvZ3fkXYYjSn0tjSX9/9IWR4/BQja0d7qHELdsYZFl0QDVoH8PsA0/oJNgUxtVUpr
xx0S9cvAptBe71CUNdUIDkMp7aWu45OpaItBaVQOTLBz72r5BGDKgN2Bt0JpbHHrMjMNjqeLWerH
WOS8hhZvZEVbbARsSnZtCBJYXn9dE/5tsVv7Kl5lcX/kdKtzFx3NQFUrVn/lclesl7pe7cgIrn7b
+yx4UC9QcuwK7s+6Z6MRt7OJRVKAbAeP3fuwOnLSBwnf5miqBFvZ2P00icg08hhsg9shsyhxzhdt
h+YHTbNidFJ5PtNjTnlBg+eexj2t9lo6zmpxyyQ1BQbdOmwuNKBiHkXy+9Qh2CYTDERdsCXoKP/Q
1WcqXj0rPBWCgXO/4pSzq0eyODi9pA5/U3WWBiAbCBDachU6pW5plNptgDyoNjlOfFaj4esPpVtK
H84xamzpZ1BIzE1KPIgTE+c6OApGO1YljhXb0gOpktf/27xJOyzCoyW3dnz6pn89n46KxqIi6KB0
pKNNliw1ewWDMd0Ytd5lRP/E2Ct1crzqPjwGdcjBgU2tXVHyxCkZSL9WsSSrK1Tt1r97WN5vehUN
0qivb5RKEJjnU552Hr1UVjgb0Ya1m/SlcqY4+vlHtW99pdDFjmLM0jWWlWSG44aPJcS2dSQFcYGk
IZ6DmhMcWGF1KXHJj+UJG5Hb0DyZ0aFnY1W+wAiFm7ftssIO/BpKHBKFpg2sAyxNqyPh295urba5
dWoWIBLXxLxMvGTiZhubfmCXvxSR6CnXNltrpaASa9kkgWjRhgYaOvhHdIswmxUQxIE1CAx86jhH
Vuv9Lfr83scasJr/drhfoi95YWE7ZeCRLY8+lAKZR0vzdKmIChUZpvGvmWayyxRCRs1YgGT1CEPw
0QWwfBb0qRoapVacrtI0N8DpcGrz6ZtLN1cVbD1XYZT4oRsnVvCKLu4atAetePb3TFqc6WQXvRDu
0ZLL3pX8r1sR2VCL4KThUGjDry9nXGVxlHngKDALlXBsuIJu4Z9Dpgi1BjpT5k9ffHdq81w+bDZ7
tzQKjyiRThEjCiWYXAqWWHXElcmYDVRG62Hv0NlyNZpF6HlMXj0Sl3yZ0wx/VMdxWWnl8RVvGXY9
KAOcI394sH+tXUScdDtzIBhJ/EFHb41ziovdIhpZ4QFKZVgZYVh4E7j0O3XpuTLHNoSoVEzUDtMO
tE4SgQS8tYnCKoyGukFKIJENP2QCgevfEeMZUHb55U2dwguU1vcpNzfXEFhwCUTuCn2UMavjjPA5
NgUDZB/lJZe8gkUY9ZM6NXqH4QVXeRi9Fz3K0VYiMFz6Tav2Bs1MMq8wIl274qf4IVt52bxxaWFw
vfIpiwiVi+rOFoxK/hKIcS3G9cScdiLiwumBrsulZlfkbNLZq43jHjqYt/vAPkwmncCYWAqSEyqH
tEAouNM25wX59nsLkaI2grELlgqyIXWapdzemjmA3DEFBkQvQLpJvMTzTn8Gwi8pdYazfS4Vw4iI
cgRD7BjBXW0B75gFgE5XhNf4Z9Am6Jk/KUv6yiq8VLpTYyL769HMOTFmIKwcvTmV61gGNOmsQwSN
DUiCyoSJknhKkpIA45EDwQeG9gOcEeK673ieKyDfDl+zqZQcZsosjEo4NUvsXZoGF1iQZBJe+wMW
8k6QniSdiJzOc92VzyiH2dI9jTklipHq7GD7fR+chiQfXr2bvNCOTtWSU9XDRYnHObCkas7+DGJr
b0R1kpNW1jDxwsdSsYqcNQEeyYYzOy76LtwLj7pp3Y7SRbIs4haRsPuj4IBxousQ8x4jr9fP+drr
lyWl3r8w1yNtECQ6HDz2TOPzpYDBWl1hC2/nj0GvoPvcVa+lVIhe1EYWnnv0n/k4ZUS/xqTM84+r
pwrG0V8pETX1c++ls0xhsERccxOZe6f/kSj75KWHzuEbkp3OBE9Zi8/HgbUlaF6x6iJSt2NELG1g
wYYnif1tJQtZ78hwXjlJzAVwlOhQJU1PGwEB6+1sCoX6KT2f0hbqBmMzW5wdvOX7iB4v9QBUUv0y
p2joP7KsCSzuDWYulV4Q+xFfCPHugZwjzq8sKqh0eofWtyU8/JxmpVqyj5H4HDcV1RjLe4yCtS0K
CvJOneDiQVHlYCj6BisEe7sLGIIhY1t/ZwhaUt9xKRtQVDtE5gDF8RUMaa3xgb4u/5XpfnX9wDsT
hV0MF0JlPxfgT2HZYX85Zr0Yhs6n7SsWmYiY6nrPj/WVOPr4SW+vey3v3jaTqpaLNl/q+y7EA+Pb
Y6htJeixpfCDscDyhakmt5GN6VT2QI6rqjhl6Ccxm3CGrTiksaGc35sAq5dgJ8ST8DpHSHtiIUDV
EBtsYyt3K9yrzsuN5+UnqCgrI7Y/6ZfPU62fc54eLBLvRkXXVUnuhBdb1V4dLS5LEIu+zYKrY+oj
Wgfb7oiqhUjfxKmeWZT6KC9apYyFVINVpD/W7Ik9787Yr09jboI1H4wplbABRN9X+sRfIKGCipc9
773J0AYJuDAMaB3gUYAW2QfQFFUSEJcVI1gfa6LDLUAJzneaMivN3hZY+InEQkPdqiRFIsaDvLDD
WKCNNSSlWR9qcwZzoxZjp4wjbsF11P2/WRgHYAXTJm82FghzGpOZK0gGDptzMFfdqTSpaIeFmIzt
2fd+Ka6FyQU84nwkumqDwsQL4fT5AwGGxFSJnEs8gkS69UjHg9lx4ISVm+xupfMhM2hOzjnH4weo
4DQEe850TkNF41ee71AwjI3hMEqHLwIVlka+HXV1YfbJMMH6tqMRlspWnAjNarDaBXbik2Mlah+H
bdDUbL3AiWGechYYURn8/9K+xoI7SOzVlgu7U8uVyqzPpBKgOlwStNKXbaGnfu/ewvGAMA6ZAiU4
60/PixCs7Nlqhr0hYw4GUYTv+Hn7ty/5eY10KEOw5l5Oo16qMH/0JPmYeIOU+9VOvHpqQvQWyC3z
HF5hgyhDkkqrE18ZYaT2kAscYoEK0NfnMleqxRMx9rMaDny+B2SLvvtKezUbcDlyLY5C+a3SQ9A7
UZKQU4edVKJCgLPxK0CvFOt26/CX+74/AMC3mvvo+Nn3uk6fWP0ZjcFSZrjjSBcuRUPVj2MPW76H
JW7mfIy+5zBZ2k/v5F+Uh4dG2hUpz91K2RM80WoOyMZnqDKDPVXowwXs5Q6dTsRemfjC/yWhHDm0
OBztoFfFjVpkRMU9whraTCpn8iPHrz2Q2I7itgux62kLpWgSsdkFMC94aR7D7bqqrM9K+nFS1jV4
z8rhMQ2lRFUXO9V2mx1dAQ+DzKu8811DFBNyPzkV4qm4jNorh/PJl7lWChSVe3Oz0HqB+qQXPpdY
xEMsj+tfPt+yjDama6y8+q+yl0aNr8txar9UeSQOc2IImCbtoGwdzwxLPVtdB3cnqRsqwcpfBmh6
Z5FDzWiyjUZiqDU1I96+xzkD7VyzuWAAiBRpAhbdt5+l9FCC5JNANHR5PhbPcZIpIu0LXzFthBFu
Gf04G6H8yHvzc1KYugpBB7KVo3cpuyrPIzbNWDZmrWDkny/XnKpBEhOTSRoUC6hZ6VaAVekfG9H0
8NYPo/rx5uWhiO5IFSxFl1bF5bKvAMpRsnBMSWFfPySS+A6ntlBLgyvKQj5tpgmmAZANXPfF1a5y
WAmk12ERBKpO52KNsJQbBcrox1NqsKpzmXlWW/O4oi1Re0i396ntkMINfO33t5HTNBmKAEjqQpN/
k1wBs5itYpQVu2p3yunZ0XuoNmPWJLU240+zPqvlV+E6PlqapytN3jcCeMORiYILR5SoSbWSOkY2
5JQtW7jgiadAdjqtWwSQqdWu9jPfbotkssAZtuR78h75oClvYWv3eTlFzKxaITOd+iHE3Z7hfltW
rSK35ZRpWf72uqSWdowFxNa90ImZxUhyxwGWb6W3TP5mv9gQs4Ay4WhJoMX4CZWdsylw2BucAsB8
xIZ/qo4gmK8XOwjznKDl3jlhX7Hwfk91AzXVg8uwowqiDRoH/rUVrMmbQC9lZcLkTgrM4nBx1xoa
bZxCPs7f8xHtsvvOHuko/NVG+r3KHjlZVYFIuTE2eAddzYsd3b4vMqW30AlUYIOrGeIeQRDpxOqd
9o5CgQg5/jt+4YBJ5p4CxfqS3Z+9TXeBEMqvtxiqZXzbiWu2T+AhlF3ouvT4fJpUvd0cbi5tOHPf
YK2H62PgMxB/+BTWSwbOKa4K9xpnHowDMnaO7D75n3NhiBLAwo1lNy9+riaOmGi2ARBAr7XZGCsq
c7+9fryzDFJ1baMneSiOFcbtS/g0btt8vRtw5Y4RPC4eb39IcRaTcAYfuKf7Se6jVKdfFDO5+mxr
RLJ3cj+yw36izRwx6B+6czYyzxq/RybWL+We4DqySVWS4sOgzuP1Yg/81CvEPqTx0v7s0O7EMELU
obQOKkbxTbe3kmZ2KenUemZvg/pDF/4USR5RqkPOGBwlylukYx9DJTfzAffhmNOPmsQdc+3XiPdu
tomJSbXDz60qx1fjT5/sx+3otZp5NWnarH7DbzJJb4dQAOG4kxlKgl+08Twjh3gcq4KCXh5VqUlZ
U8GOHWjtt1SNPnqNbokaOFI+/rxg3VsC3MBabM30s2miKwf4/cvr9gSycQqeZVp+t/sOvV9sBGdL
wQmIcWolIU7GbVeTpMb0CtOGvDBFCd436kE7ZUaXDR/Cdz0KYm0x7pfXXzyFqjdffKEpPaxmg1uL
HnYki7FtKP4+wrHMR1xAvtLHj3nphQflpmmLKde8HON12YTOoft6AJ/FiztOQux5HUaRnQqlmyLT
6aCCkXgVcUSQ0dukHjPNvAe+oz3jf+gGJWBG8WCSX1WOVnTk92a1/lt4AsRT3Yb7oV2h8s25ibL3
ry2uD+yS2xRIkJ+tj++OO567SXs8GOgRDnhiGJPrfs5RdlJW1wHCFuy8sdKo5mGz8VVX+h3CcaF9
tAhO+0Dg1cNDYK8B3ircrhh6wSqPgb2LPNjT/W0026yNLeD+s3tYxuzK0pE9QhiQhJ5i/SUh5Jl+
nIZSlWCVc5YFv7qxNXeGyViGCS7J4GlDZWLEpTPJzZrr1pAbMJwAUVbiEq7N5dGmhTk4SZcMNFnj
S5HSk4hHiNx7coUFEDmFT5gx9FJNR+M1CyGGds03I0EvsH5Ys/SxDZnwVSLEKvb9BFyUHxDMARzn
t6LWFaWmIlhjr7w+O0hpfrzbhozM1CUs5IzrkhlnTG0RqDt0bCZbUfemfZzwPREDEz77aAKD4Blj
Hc8Jw1d3c2GFILg6K5Ftq+5WSHzr0BagaHok/hLiKKm9E6nsBTC8zJg+q96ZxiUJIlKmwCG4yPMA
gwttnu6OsrKkMgSweHDzRrNNr81Gfysx6B0ZA5odYxLTEvQUGPHv3q/l/B4vsOofeI/DkeVApCfX
qQ6fOgu7JaeJfDtDopKyjxDdBC2hYtHqSb6+c6EZp18OwHZOAfD43y5EMR6gQ6TdrdCG6qdykfr5
0Zx2wvQUELHSqc10JsQjd283Gk8pjO5y/MEnfnemSg6du0u8r9ufCV7r5HNefMvsFiTSIh6wlhdX
k+FSJWw6hrBICFv4ZmMkoZdkIYUsMeHKhZCSDv+iY0iunSn0FGHL1Lp17pFCmI12zyL+ECoGUdj9
ZStoqkHcrq74WwhfwJrKfoZWTz0Gw1xFO/h7TfM6B6hVq5X73bZtu0gfLRuNsrGvdxqMRfTiHPJx
orXxbbtoXWln71xqX2ziXgfGAfo8csxN/qu3VsoTefUtMGexMA2CItiy1vlsLeYglW3VVEMbMkZH
Og5ZlYNiaiFILjMUH7tDxcpI5+4BiDHtlCbWQCUC6Tt5tIKHlVjtuduvUfLAEUDfsMQJ/oXxPj2i
Ead2yA2sp5QT26vu00/X7H3o+Oizk7E+WZlhnzgs6UYcNCv6Rv/9IYqrXaQTiz6r2nZzBsEHulo4
vYPtxzx/As/VX9cJ7b8oFXyHv08iGWGLHReNfpC03kGyNBzQbfl3LqvTHrn+/flfyZBRcyShH5n0
HO67CmLSTa4wpbQDGjTVNnA6PzEAqDlwun5iZSPLjEkkepX9ZchZ6l2IamaLywj01Z0PvfsvlJUE
YT08bd03AU/KshtM9sqDhjj4XT9cpgNEA9CitNiaYWBI07M7Vt/sdTQoL/z4w+JSQz72VVK5gcKG
/4adaThQC4bYG8S5a7vjVKtsOfS7AHaRW2UvW1WpoWa23vrza540Pb8kbCPGVPwLA7jt4iEkbAjr
35mDQ32J1VpOKRJHUcnRt0e0rfgXaewAzfqnHlb6m6EVCBMoTF0GqOdH4IvuYIZDjVyGaaefWDcF
jhrrh00E2HgFx0cFzEgCTwls+iVnuJ9gpzTCavxcTqE3y4hoUw02fQjI4p5nZ8HNH66Riq3ZriZv
fp2fI30tFsOJHi+8oA5q9q3jCEpwnJNslbMcCwww2SXEcthMoTnLXPFzlb1EwLnomgczoiWYQJmE
AvS3W7VRmxWp1KflX5uffkThTC/1jr0zvM9NfCPhtYqT3g5G7JaQOvNTLn09vV07jDRNuy26KUNJ
5LbYAh352zke7u3Xx5JyZxUreo5vv+ub8guAQm1XrgrXUagi3K5Cm5Wkn+5gmSXHIEmmiEjtgH/G
nNTUUP0Qhn6pH+1HPA+ACauisOjPFGJlIBozzZctRVCT6jQXvWLbCSfGaQfF+aDTOzj/zYCw77Nf
Clu/10NwKD1ju+bcKOD44jaDLyrmDtXah5HfReW42A8l05IPT/uwZT2gItLA3EarVeaV8SIf8mko
o9YS7vXPSYUth5G3nyQRNr6gY9el7UI/4Rw5KEu0trtW4AjZEsiLKIS9aU/CLPf3Oqu9qZy/zNog
3cpF1srb2D3zUnRsInNKuhuqaQFxJX436ntRjZScLbdqmoPlMySodUEn0I2l5rWeySrzEJudAOfn
V/GuAtuO9qRiPjhbXSWTwO7VezsBjWywjw9LLjR7xhALWzoDHAPd+BwB4MYR6oPvOkZRWHCB/RXw
Wq6I520crUd5E/exsXZsyfHv9FEzQZhVRXPfXEsSl5gX5eEBUezSb5B2PGSQnLH/eGVhTgdVBOic
d3dIMiVaqe/A58YlOn+DWQPMThGrRhrJS2qsb7d0xVkdD133RYVveEHdV7cZGV2gD0b8zAcghYUi
f2EJa+0YOG1zaYCT8hkLQwos378X1x9s/WDC1QClNKsYz2jgnMhYJVugK9B/hAhrznIciYW3VP9I
CU1m9QYqiWxneaVmBTLg8X4OO134UA5Cn35iryzyrxKCLDlYAzqH32lro3D3a5g4fOH6H3RIKOw0
GaVaFf6lchw5X3fOmHjRdaWqiYvG610JY4VHWgEEDJn4fqTEHkFAy/4dwF6kuQcHSlc1K8fNtOee
U0lAtoSEDY/zHlp9MHlPTfzjBI+rl7qtePy/KOSEuZEqS1yKmXJuuUePVGuA3Z1dZDgUMPH+aPiH
BTpKrqY+dHoV37Ah7oCHXpjWtcYxJdgh3wfBUl2bHOjUFgWAnJcndNem2JOIHKb74X8XubyCyXUe
FKkQHIPvJTKAGMMR/T74c9LO4jxH1xpEZgLHt0zc9QSKMZrSxt/1qYxVcJxCtEhqLYiCVcY2sXOM
Q8GApde5TGX+HCIxYm4GZ8uIDIfUKMeW9H2Nl0SZ2lW0C3JXDkXVJVbdoR3CPB9RWqvlQeQ5MFQC
avN8ZUtoVblBoIdXfPYMmnNR45RehqiuGY4Dz4Gfq3CZpF7XUtpVnSCYTm2PmpC+bD1dPvVXWT/l
L7KXX/rf1d4DQTiyB0kNqYLOOXsaWEjU0sVBDDA16NoNoXTNhxGPEAua3TPVqufMHEz8q8tgFIUL
6UfBj4zIz5Sbv3ghayylFA2s/ySgSDmwWBZEfznQ1vfc/daAgF4FNiXAQM/wcfLxqyrYYUIl1L6H
AnOHL4wG837P88PYjK42BytjjRWdlshbiT03bECP/Ne7fwmhiPTrYEvHGEpwyoCq1AtSKfVHWaYs
UQOddVd7GBQxhIff9zaFWMGll1k5UdG7PadBnJGUBXduyiwsV3XilSiyb4zwadIrF/BwYT7rtkY1
jT4mKv707Og5hbnHzYxIUTbRutd9NkgzQaQDu9/qYCQPt1DqYAGw1Qe4YkhNOpBXBXF5vzFFkzYy
qxx3I8fR9WXnCvKyptxhj6S7u+YWHZFy1sQQQAS7R+kvdtSePmXv0Czf7zoObrjXXlebtXL7wR5G
1uXpq+ijsHzVFFSf4otHQXm3oTsVkWVmO8bqfEdsc96amsSmFP50K+V8yxZ19pvx6MGvrJAcDWEO
MVEfhuAKn7ZkdZZEyynbC2YiIH/xpA+y5pMeGPUt+dGryHJmcZ46d4f+I51OOBgLtOIkebLxxGxJ
bIj7Z5aSCnKbEvNKJd/IB2S8MXw3Q2BuT3xYE3jggQQDkfclyqSsYBvXn43mp6nuBkH1xXu5qu/f
6f3DsE7RIHUtWnE3izqkMygJU+0uzRVUNI9ULlueuEJfNOs9FnapQlbbOr2lxcgPNz2LAbgS3Q6O
Qa6Ppa8t3mkjlrnnlTJ/qaRYosIc20E9UohECJZj0HOl3nStbLhLgG3I6X6kaxAe3HDgI1WfTtxp
AGlBhlKy7aALJGu544gFPf+lf7TJjsXaJzUQeoSyjkhICpOSLn4RqSi2Vx1Zvood678Z2ptF+SV/
xOpGUYL6urlaA2lNuHiWvwLMAYwUwCDfBW9ahdtOcPac3fhlVivhzYWk1MQdkRMBFVqsIjoRuT/r
Ia0/EFG/Hp5xCE9aaBfQYeO/jAJD1yjwGj1I6b+ETjPXbJeoCokVd3A6cQV16M340mQtNbKW8Ro8
dME0eycKB2TuxRPDD9stZ5u8eJkrbAxafMB21l9wH1619ZP30UVxcDaXI7Z7vKSO7nSYsuqRzcrF
6ZdMj5eskxY50uRSV1jkWPJeIHifZk008fzMxC42pEKZgDK9qPdUon+6URRqAAcujqLctxDioSfT
OWtwvsrH3VTA2rHl711usSoJYrmDXjBvMA2dHfeeBHYkG+Io3RsV+pgwZrQELrOKaG+BNefzzk1E
xNDxT1sd5/qDTropmMcLLC+YU39zW7XdtYDlQvrKMvpjx25s7rtq+dxhenNXSUfZy/2PYr8AA+gL
RDi7Qm955IWY1dJadIU9CF7IfoOMm4jZwocxTDaDitaper6uw033OmBsCERS+T9H/kmD1N/2dH7b
QZk56QIBE9pkY8XzrZ+qoPMxpYtvaKRXJv7HWN3ly5dvd7OvX8Oi1+ARo46LCVqPdQWkQwHyLrjc
u45sUKxTqcS58uFlcj+dbIsTxnKhTguAqh2ZFxEYuhpAyb90JWuuVNCBzdTiD7176g8Uj7Uvu+yn
GxMPZHE96zuZ1rXHZSX9SdUa2Sp52OfJObkDoFcRepXBcMhAE7FW3kUUzQup+/9GOgqtdD2vUHyB
47pdtMKEr/dQk0S6UZUKTaFYmiFcYprlTWxvV2tBHV19nwJjt/I2g70glQ8GTKcl1rX+MgKOVBb/
6TcCH5e3GVApQ21XltzZEa3tM4o079I+YMzVuagmq1uCLiG3Ml1MUm881LcGy8rXFCkcpF2dA9o9
BKE3gnp4nd23eLacfzfhA8dR6kPswblfXhJbQhvyJEIwYmxd/BpBTcHvBRhYF7j1W3jz68J3KNIz
Sciv0etWjosfOsdWO2T41sL8DRkZ+OpDPCld5ZblTEpFF6NRlDFyxVTya6Rwi0uYPplLjvQfr/Lb
hRBoymXjipdfL0THCXU5Af2tB9HUDd95sq56Jsf+A93sFTRxV5hSxUW0/jsu7oHJOXzGXto6TsP6
qw2bw4Teal/LNprqzyAjs2IQchOSJgir2nakG/V9x7tVKOjKu3iZSLmLR5wdpnl8MSLhWNvnVsNW
j70QtYPnf1n8QkMmnfPG35O0KeXboBkd6dRgwig1Y7ULppNwaRdtDZ44yLznYrCM+CpvJDG/eQys
FgZJaEc5ET1PXnhdFQ4K1KR1RZ74TbyFe41+5dh2mnMkbDe6gkOSMtczg3nJnZwe07v1FbYmNT2l
FYsgQuwVse+a81fQz5Hi1pjGElDiwKCsLGHd9vMP+gYoxZvFLD4eLaB5MR72huPGNQT5mz9eYoM5
VX75Ba35W9rNXEucHeAn15iQHgMdsP6ryxZJ4uhZK/o5DI5oeOYUY2LLBLCJd9eMx3MzuJeTODWD
FI4ag7brK00Nmn2+B6TY5l5Wv6hvRBTOaGj5qadUDEZeJX0fv6tJbERktvpCJyd/Hv9K99f3sUy9
Mf21TkSwUG7zZUMuAIMfwCmfJoTyxXOly6FF61CVUckmisF/oQ2L0FFeU95kCdDN/H1avx/OYP5v
60VpVATv8O6PRhZ9BWHFLDQY+Db5CYJF8KsFqi58xvY3mTc80XTca7gudJQAL5LMlfCqsefko92J
fJNgF+qk+8d/X7whrCKEITF/XHuXrObWEyilhoSWAl4ELkaiwaTpb7ZkExmXXMVdeQNYMW9DOitZ
He91rhSKDSWsuHLWMxEQep9oMcAj95puY/45DOv8r8dCQ38VXzsHGph3JiIhBbsf54PfJl/s5M1B
S6hcImhMLtcYdVu6XWUs5BpW+vEN1vYODVrjz277r5Jt8X4BVxVEByAFmbCg1kuOwBMtrJIEuNVJ
grd1KXplwu5wmflr6+2zSq3F9X9KOZVOJs5ZKCe4Y4KSbxgMzZz1KDGl5tqoFG7m6fKvPuF2j9Eq
rGSzJQEkUdBRRuRxASY7d+chZb5TuNO6LDqF+EbEn35p3UwU28YvidAsE9bl/ZZOa8ZA1WgE419a
TCR31ctDK0LgY2ZP0uzf2BnEyenlPktA+46ErDm6stfZtN9Ts2zle3aOIIwrhnv5TPx7YFIDPTjO
SSDmd+J53bc2AogqQSQ8j8GSWjfyviTgcKc3iqIRdo4LfBJLvSduQujwd4jZ0g4oAoTGrx0dbrr1
ZufeopqkLZHEMvjqjgKGZJ9CkWlZADOVyWxTFm1jgPd8jhSuVvafSfPWlSZR5oxLBbrbQC2BNj2b
1oHeHvBdL0Bx5sJmWtOJn3dTTHq5kOdZyk6uy+SXKLHp/pyc7eEBqO2RMkg/3kY/svIpRfzfBlRR
wqKWuy6e5KIjwOPFHGSnISIBiJUtQFAvKAbofnt8t9JL5sbOtTzVl/BSRRoLAmqO8vQHOVG3CoLh
n/54NVePWxH/F6QCjVNeutOUAFNVvaaG9Tvp4jIceKNT3kTp7qbLEcbk0fp0ImvR/WpMm3yKq0wg
UVGGnlHbOzW6b1p4sCE5tb3SZSNsvbNpHGqfio/cXHnrWhn90KttWUjJzs37F7Q/UGEG9MwiogMF
NaKsiDOS9DpDBHZg9CuXn9GOBfTmhWavyFuDz37pR3Iz8lQYmfPUhw+fcf3urtSb05pB9NyYIGN8
i03ulqCv4t/G+wZURK3c4Y0kE++ykoXoeEXjYPOEDZsleaiGSs3Ga1L1HPaQlHtDa8zQu6jnmaEV
KgtpyBpP8ENhBRyjmcfpDnWtNWsrJoqaW7yPe4H7COTD67tLYuoHH9VT94qwSbL0oRtSAPQ9J6vB
52zUC0L++9LXKVwUuHGrtnoSs1tszK/UOGKvw5fhmilLytOPd/Tnxex/UdsJGnW6VGtNt/bDvtET
okgGNL2sXJCzMPNnxlGgL+r4FHfavdW3j1eiwqfcb9doBxCdARRPEeE8Du7w0obr/bzZomuvS/mx
Q8dm+vr7QeZD8wfzeT3Kg4jC0Rio/ndKN6hZaBazLcak56hbglPBiRASbo+HUZ1XY/cqDCtQg2b5
rN8R2VuhOZ1VDW4iEeROba/PeNrdHR0y81Jr5SEU22S2Vh5SigQ1sF1VepEJCZbmavFDjABwqPPA
igB1/c8IINFX0/R4NcZm8CCHbRB250kMb6abwxaqQbvFmntqtJTnugv5yJVfS7simebJ2pO7kz2H
qPicl42Tl7vcGAtMmTMiOh0uYXwPUxnInxxMQBrLSCjDHHj9YyV88wS4RZl7g0uuxAn7wv1Vll6q
2S9T+I80Lhlq2tEhNK/KJgj20UyagXonKwmLYkBdwkRTwoqUOW+snHO+Cu41MslVK7JDtcpkk2FH
OxI0oTFCeTSKE52Gr1/89Bmw7191oWtlPxXDjCvuO96N6Oa2bnmCbIw+x334qN/bOI+yQGCSZ8mr
7lRxcbjcSWM9T5a/31zsQrRMYqAovZdUmc4rFOI2m3f4ccEy1OqdIGDT+IJ9upQvvDBKpMi4QZ+/
Q1NzOTCm8iuR9gFCrGcc6+AB0GrrrIYXaoAaTBUuD4lX6DfnZ1uQl+QMLQV7HxZXZR1v10HyTeiF
cyaXRS71y7fCy/sL3IfoLEhMfhQHko+r6qsnSa9/rWeR8OvI2a1Kzci9sNCZ6d+Q/hVq4NqAUj1i
jShKvh6dzGvAXom3D/rBzVBynSyYunkA4ar4PDJ83vM+o6nTuhG0XWv5VE5yJT7mRBA0ALN/23Yc
YSf2QKqVefgFGo3NJ+pXA6mcIFesRzaqXE7zueTMfOZy750wahSAWpOnHHsFcZkYM4MjDJaNCeal
UK6R05gScruLsoXyKfKp5YPb3BUVo6ywxhL1t1rYainHmubq3OzCnZ05dzvUKjbAeMpapERrWauO
gJQ6TbIkmILMK+0mddocrhw91L7YboYSjNXiInTmOWfI85U/vYLzKbIxQEo2lSA/ExTuXIXrs06Q
tFVigw/swVc8kN3jiTTEuZn1w0v9Ka4R6E432ml7u+4erN880HNMf+sYOCsn0HXwL83hVcuXgI0s
UeOO1MGl+QfP/yn8KnaPrTxiip+DohcD/YUyDIBwmWdhqXee2vQxv32THhPIJpUJPDOqyUsSufzd
Gw0IF+UobPotpFC7QCPAXKujlQ+PzaLZ7kF9PTBQj9kEQLaD/yVSbD8PqCw4GGVI4cKMc6yImJiA
lppkDk1Z0J5VE1tlIR9Dh0pzKm4rT2186NlCjDfz9l6JHNbE65+tE2ozAJ6PrjLtZX+Xxdd1lcD3
NkjFj2xaiCH4xrgNeCZnRmc/7DKHV1ats1pz7txy/Y9E2jP2BMg0NL6Erolbe+H1NtUnLcC5u4Q6
TwaacyqEu9shd5bOI+qx+09iDpyNyyi4uyjcF3MONuPKRR/g0AekSddB7iWaiqH/+SydqljxqCG3
H5Qt04zekhI7kjqOxj2bMr/zCAE6EhkT7CrYP+dneWYOp5WJBVRw4hITLct8XPGRGN589Kn26d4v
b10iv1/5rVmQRc/RP9ZcN7F1ueDpWL+Hsnxw+KAWcquGJqDJZF0Dya2pHAv8q2Z0KcAurXq4FTk8
7eMEonR1ptQFIjUrSubwDkyVA3+tWR/DZX+STqtm0Sb0MR0GomsTVglnOWAmi5rJwEWihY/qJnCm
ZOtJiXn/uuHpl8+2mC72FBdog6MBhfHDbug8rDYTg+84jMEXKSZ38ma6FdjvoCSeDRThxNUhNB9D
M5Ec80eXhr0QxPSdjtxzJMCYoGI8aa3sfqsyk0XfAJhBiFbn5bkB+ZE0hq0RpzEA7TOCcSE0EJnT
yoz+NVVVy+p+EAcxudUa8Btkv+61owMbmtlFtDVZly4Ka5ujniVKjOaqwbTnSahobfnxKM4AKy2R
B1wcyJKbmMzEKLLMz3C36WN6Pw39u9gcOzyrFGkrfP0KO3XuAwkGfTF24CX55CFfuvkGaSRdgvff
PmcJtCew0xYwU0dF0/0G5tVJj7ebSkrSZkBQcm4zPobt9e3I0ZNFBTn3Z9xUSiz0fyQch/LXG+PI
yqh/THFlkPBONdM+y3bD6biXxHyeORztccHBOCf+7YcDdp2CXxbZsZRwRTPX7EkgRnX19//4aS+9
m1TWPpCqR7uBZf9PNasGaJlbxUeUl5mZfLVAQkmlweFmyktswsKbummTCyCu/yGhSo5alW7BHfv4
51xhXMlGH8Co/XVrqw4opUSUgEFqQPZlANQb0c0+srYID9gDX55QEE/3KgsBKygTCj+VKv386r5X
cXce8FpXwvj9bhYdKvZj4UhICZT/9EzP0Ik7ZkQR6xerKnlxkVqprob4mqfQKSiBDWVBfLaTQefa
PJ/IALZpOK/sgrEbdH3ZCP2lwvFtuP4zh4bSStNL5iI3t0JHra8slwye7EsrHHAnM6bU8mc14Z7w
nmSu3uJPlWKFu8WR903ioDDTWr4jv2V6xweDMH7eB9rwOgo77AmQS2NvfXLrgplUpxWCW1WuC/MM
hxY4g/gf+BqTz/ZO/DAcm09dIh4mg2ywKkwe9OYp2yEpmZmAY5CNeEBDpqZDRGWv0IXsgsrGXVd4
diufwygqYc12LSiENIkNfsLpNy3j0pj6krcIvL93KJmSjubjBycUxkd36LrwNJtFex/qy0Xk7/L6
LvgyGpbuVZSUZMDuXHpAcHj7H1ObeFoPjd9FFyHO6XxcQ+4r6xR36EKOWzjreo1yoMGGxs513sUk
pC5PtWeCbhMuY402gJlPUD2ncXHWQUGKBpupZY5YquKAq0aJZrR064o3VevpWvXI6dJmKl6Li40t
IRBn9LN+Dh2Rh7GZZPV4AVHdPScvqwlSHqGHCI4fmNW9w22AxPaUAzVGKISfREK12W6/GaWB5R9t
mjHfilGOi5A15T65ceSQ1xmF34uXayotqkPor1TrvGu/fVBsz/n/TX0txA51oN2v8ZOcqelijJX2
B88leO5ebgK9qfum7DpF6TlHpmt5mHzgXrME7PXrtRlF0Ie01EVUW54T+DXxnMMaQTNiC3jNij0c
EWCa7uiQT18MyccY3P6Im3rNP1cbmz3h0bhOE1ljp5uZANg7Rw/uv7DJ0EjMBVmeTtg1G4hpRcdZ
lMi2tQObiEJ9DSip+z8BbYvmvlBqkDDjQ/oNWqxmvC5cTu1y4rI+3cOowJVRi5FxtT731EtDtKo4
GcFEzm7XQe8fnRm0xGIcr3qUArlSZ7ieZ6a2QhAay5dFN9bIydGuPfaMXDFGCvpt3AIM/Ss7CagH
qeU/wzmGFxPDHTF1FHExrUDoAVXr+DIoDUwZ4tocGrcikigygl8IjcuwOaZex8YJ4HXpfGJcAvBV
W5mG2SPMN6oYdtZqRs6bdGQUFTDjmywo4xv0SvonizDPKkh+mcc5bdcy8O088TvvJVFpyD7pIxD8
K7xheYfXGY710n3Wb4oA4gfrMOLZhC/HpYyoZ0bifxxANZDhv8kgr4wiT7R1H2qyyaKMvTf02RAp
/dFnIkHbjiAHuAsV1domZSxGjgRsNqQCl83xcDldaHahnSE8JJYFU079kcSB7/cbJoOo92DUrkiV
NjDocN7XB9Ep6UIS8lmS9hjqs94mOCmAggz559V4fuUIMdOCoOFJVUEb1zuectaLb1MMa3zrsZ+4
0W+wTf2Mare/n32mF12vc0xDxGGfCtsZ8nVWntp37/XTfRGSTvObQlgq3kkVHY5P1bXo3SK911Pz
vogKHO6G9DCBuIbb1lTBAnRREgj7jDHgLPMoZfJ+GeA1+G3ThY2toHIfgLcQJk2i+OB3llvWonin
MlDKX5SDVcj+KrFgtbVmW3jq6Z5yaeJoXHmxlemA/tccnR+xT/jarzGQ0irVlg8cfAVHMJwCAvu+
kw9YHnAQt0Ig2/sa+00yJEnls5ez/NOjTjBqsDi7SFPha30B+3fQLTpcZUgENFg2nUgcCEBwITc2
pUQarEGjkmy+K2MDcQYhEqad7wykmzt0m4o9zMr5GyqXtsfLcCmNQjS46NMgpGFcFEzDc93nifQJ
ymfP+BlUw3Jysfz1KbiE8ApwVKdKwBYyfFHIjWoIVAoTOLqt8z5kb/c6lmssCXBoAbyNgA1n7OJ5
dfljXaCqqOeKnlaIxsB14/w3jXYr31rKfTamJTiKyNqxr9Pkax70usz4R6aFXSxziG0gqgfdKyot
QFoJzq8qz7zpGQbFXxxhaBj8XqCYiX4Txi+0bEFbuk9iKWD5FhsuhiOZ+a3o8Qq+4JvuFshanRN3
L1yHO1BGVp1R6qABv+Ic19C6vf1Fdk8EduVRkJi5ESNQ71TYKmo/IPjpj4Y/EWeCl3bMak/bGXCH
yjXH9SxnLCa3gVKQTCGxeIPbv6Cfwhh90n9sujDUXUK1q43PkJjWBuABoG1gefFZcP0GbqNSQTCY
yIbGFa4SWVk3aEuPwtlQiHZ/JfptRQW5tP+W3fKpMe/VY4PIrlbsYuQW7oXDd04gkfEEnossdU83
N81kzRbRTZqWlyqkqe4QUfvAhsfcPQelv/9+LRSHvbPXOJGLoODLkhIXAqDo9Y3F/Bk1jdZKu+Jg
8krkFvZct8mHu9gFzXZvuphngD1FPx7mz4kuwGqaatj5yy8Rl4vhp0/J6xXZzfulJaA/B13rYkGo
n0nH1gD429nY+2ok/aGuIfqLPCYUnskZDg463xnrdiTVypi8vHH7clBS3NMUmtb9PlsaadcjVYsh
fOK2SWBOUMJNoKbRGk5w1HiilbnlUwBMUcCW7CPlgA5eXCNXJM7Qay34V4Izme+P9uop+O25rSyK
PjGbyS0H62LnYsL4KMwTYI9JTGyuh2lwLgH3/dhPXhWfZFfsgHYnOHIZGw/LmpnfqW/PqcLUeCm6
76GoTNXXPIe5PJwP1UyBoZ4sfLNSq0jQBfN7PDPvXcfIoIiP5qa684YeFXYBTEc/Ad/Sovr5OURn
BOUaOiCYxRLcJn2/LrYdyIaXyXypvz6DmYtIMAq0tUosKTuuSJgV862ZFBaVi82wtubrDtvM0xtW
OXynBoCVL/BGOo24JmqnF8a4vE0AVE/o+buXrNSHrQgyQhyki9F171NteRk3c+7qX9+iY/zztspG
zMs2NIGp0R0aIuutvKx29o6yvHlilz/8dPb2X2e4evl1x2h/eztdAdKf3sKAjRCcYYKL06mJAR8b
NSnXt/2tOg+YLuThABKAnQRpJDKb9tnko1pfBMmXptk+RC93v4dP5XjT9+Lj+cIJTpvR6Kljhw8w
cO52cgC4vn4TaLQCo+XKmrWOetug8RUSnmQkF5j2yi6CTTShQUBTNsJr2UoF8lk4bEAr3gICiReM
6+T/sO1VBRL2TrpFGuhcUF9GKZIuJM4s5RcER1Et+SvPArh8DR9YGMnpWl8mMH2zoWoNsLGq6zz7
3fPfCoud/aAnsZtvpYKVXOqAO5oaHFu/qPOZu2E0WixKRvbo7ps1G2Lq3mNpPX/lyGsMT9zlHVAM
SJ57vUuNHHoekiWIgLEXwAbQoOhKJ+EsReR6/fCXuRet/fLe8TeZ0j9UYIEdD+2bnj1dFb2QP2WD
hZ138YLzl2aPNrN+YK0APUbBGx7f+HhHk/BjzOLmuIfcdqnAeqycL/XIN6OxPW+A51hiQ0oG1YvG
9TC33LMbRdpsk09c3n6L2UdYa/NN5Ef39QIGysZpiMGyTvxYsY+Avpnp3tCdyrXD8G9kbvohrwbU
HmFqZD+wMTFaFzV3wXN7vz2D+5jwz420YukbjGTr/JIKacWnJyQqzDiMVDwT7h+tS1Aw4HMLwywb
2JAhQfeXD/6KGCf14McRteQXBOJ6bih8qrWGfmAYrdEcpLvntica6PX6i7hZnk9/iblEacccgs98
Qk6pB93KDyjCnsp6bRDsacUxWzuJnieh05zQvpTkg1EZHSVIi84P7fAZBaURiM+fWkkNlLpwRGUI
EQ+iKsi2Dz22N2tdK3B7V/6eSDVHrTZBPMTg4SwUBXPmwy1/xslA5lY+inxEyM5kGiUWBXcI+q1A
hgPI/YMZCCJJjbOAM2bu+tcRflJ0iVAS/cFwJSdMpz9qhzxuTcDX75mMd4Yje+lUVOmsepLebjlx
4ORAlzlYIGfsXmUUXl/q+Yub1rbOSG0Sq5dFgKzL9dfiaB34k9r6Efbf1BLybOg84i2E5/QP87bV
2iMqWfAXDHkAssJGZ6sOcfyZnEE8LmPH6h8vlOVr4xiSzll2pTZ08obGCsBByuCLrKXlE50hCn5k
j+JTxEtQ6L8hee6nlIbwnNA/2TSKSAlSiK1LvcGEPspIuw6jxJ4Ppw65LNpCPdBl1j/fWEfN5I1J
2hQ1E/ZiRDo06eAGT437ROzNPIUSVHv0q66jl/WaFyCltMjoiVq/j40ivYT1YaSclmEbuo/JzxLN
gpuWPr27vaitSqYupbUFqFBXz+6NcmxOWx4afBUp9EgCRjwvUHA4Jl8EkakwSY8NDENAcFc52hO3
e43E7l/2I5kwI+n8E7oVRbFxrpRTjEbLgbP38w2lbpY6VpJLqU4VmaHsLKipyli0U5KtwMDNByGf
klIITEYCJwYRfuloxI/61rG1xbmeJ2Wn5dzDPlOih+CzGuS6yTBIoCmn0dAGrK8V9pjYjH1MIRdq
h2YuzlO+W0ugWpZfI6GZ0uitjGmnqjwmK9L12IozjxmcOrHJhKeeW3qWgQMWmNndZkgqz52RiiVY
e31uWUvr5Dvk3uxH92EnkNP7DnjEE0REca/3Oj6VBVXRhQVo7EtgUywRyG2EYfwAoWawhDPQ+9Bs
IInpw/G9HZ9hhInCIiKQXltfV5ztn4/ow0uBESPYImRwrUAkheR/LmA142kTqjy/3fl3CNxUbYI5
RakqNNAKKkUmBIn7h+tqJuwKK5QVYh6Czd+/Vw6ksUbQARLuGQYr3dIkcF2B+R6yUoPBaFUob0vn
UE8cZwjtNeJp2aEq/hAS2zx9tTM7ptlF8crnhmyr5J5qWUeXI6mcpgfHA6oY0GGNLw40781qIoCu
kWDaTPYVga8lkglWRtN4HIKSoQGk1aV9+A42U/ZwtVJFkErfXjJyrgv/QOQXo8bxH2dnLX0Npx1/
/Ba+mZr8Zkq+2WbPczch5AqgFHyHPg2UZhcv1tVeipsVtP7V2cgS1/02crUa5o5BcUSxQ2W6rTMu
kE6PX58vP2Im1oE/cob8w4Vyp5fCXVHNjcoxfPSiWAmhFF/dAtcpsoSp3zPNE/0Vw/SPzcdwGgHr
/bqPBy9ftq70eljtwZTJezntSs3saz8MoezGOy4Lx3C8sRXqgglE7TJzYqSH9f8iOVgVT3WpLihd
51JnhHY9GoDSJiX1mX8QBpip5ccbDmnuvvnOAemdF3rOqoFpTdGPSCzSlPCwU1Lz3v7jfJo2Etf6
3YZhkM/kMqYz39mU8/YmD8hLisDQ/B72xhN6l0kSqdQxIXrgPQ1bR+u9qvZre/LFJohuMav/rGv/
NBWO3IcKsjYsr+5UPUHfsMA9aNwyrC5LDcj1WXEjVu6WhxR0hRwsd61RC0mwRnnFVfWMHnAfpLmY
vo6kN/V2Mh5tJLvwtnlLRqPkj1NYJTqjFtGuU2P7rIAZGaDgcRcWqPjAbpflfqXvQeh/cC4Rb+5H
IwBaJz+6Eq7u2S46P8bTfuL49Om0Lslu1vSO2liOknHO5Zlsae1E9Jn879uXj4HA/m4Apcdd7msu
wZjNQpvBRQwz6c77ikUQ7AomoVzri+J2Ukt6hoDTA4qIIymoUYACh72kJ+drQgMJNYuXO16/acxX
zuXF8+CIsKvWemwREKk02AA2tiHIRhJU1ntTC6TFhWsBxDeB+kfDwgxY5MWtwq8Yuu6busfCLNyA
uwToZEgPSxDD5xY5kCun2PGEU5vUQ2lx6ETQROV5P8V74Rwk91hARziNeo+xUD5FZrNXQiEG5Lo8
wmtOb9UJhRBDvy6w39w/zegxKluoUscy7u/BZKe8gK5+ntFfc2RiB2dsGdVdR+q2UPJsFg0ZLd/V
udiXEt2ePq8ZzBQtCX7k81zos7M7icRxGwgwGVvs2VBI2QGLbuUC+WSmED/e9YU+0ynIUjlmnme+
CP8sWg7P7WmW2pPh4BxI8aR2arc6rqGBwtqLKd4Tet8PQeZP/LsBTcd0SSysHexalTRVEV3p+PWZ
zErByE4WvoAO03770m1pHBUQJRaVf9MfMTTKem++Ax9iowHvlloDJisJBKiXnxq+tvwR3wh8JYaX
JVGiKLElnfJJD+ruq7SVYl3SNok0R8/+rpO7OJ3gk4NxjVRJSP4m/AAnX7bKk2nTPa/Ageg0nzt0
MpT0n0E+3N5iCF2wUqVBhScQkSb8idGH+43ifxCUX7WBXxu5GB3QZ0pAqHOMjob71xZuZ0CP/Njy
nthG0lzn4LlBGJFzpgewbOG95q0n5EyPkKau6BFpTSXl94RcO53bqgcq2iqfcm5MxZK/tU8lQsAv
X4UVbnn893ETvoxAh8uj7v3CGt+ilN9OkGNsV4Ap3jcYd8D3RCwvlKPiJF+QMJw9YO+LxPPmXic4
gy587r+Mii7Y5FuuQ4o+NaT/vkI7a7ZzOAqLZWJPG6N6vtvzcSffyAKLXpwYFa5r8oS5a6CeowVF
m3JSVeUYCyzxRw4YUZQ1ebUZs2lVmMH2zCD1VriCyATxBe10TD6HZe9uB7tMKcYWh38ytde0av9Z
U+kt34kdj3RCx0FfEDn/C89nTXTxRLbCaKnNRIjDQOpi3QKyLNa3pdvFWkb0b8c+TgkVVx4ZhPRG
Pa/CaNNjcVHYsqSiH7MoaC0XZBmMfBkavso7a4XOijR6X6sQLHRiPWsooieQoa5rYhL7vAQRTBt6
qj6vJf4UwQd13VYMIC90F8pV2UbNxQp5KEilErf11tSDxWpKB1SRcNKI03R/hBhwTPS7QzvnUM94
1mq51huDC6lvcz2uTpjgUAJkvir3IpEfTsUgMb/u8mu4Evk68v1/4HAnZtZ+7Y/wkHMftv8ZRlHe
5XrFphT3IuMCYLKJYGnh25C34OfvvFvhY0Q95hnM2YW/QSs5QiZHYldPpwpUr64fSt8I9E+C2FDx
hjlpDelNHE9SZ1KAQnbvmaCHWCp38Qq2t0/asHQhkBqLBwY9NwEUiN525a5TS1d5pvswDDcdNVT1
0wt+eSAXHQtKIXBs2QST19ESE6IwT4EqDJxaucEGM0wTd+0Nc8IcTTG26uvFUjGMxYoNE6ikcqQU
YMsN8o9z6jITj4r9fn4raTjd2S866+SnPOWn9QM8tk2lz3m2+KXXX8FNXYvVJT0AUlgkIU7r0THa
60222lN6yPffaZkTvsmAkALFLhGXMtycbAc2mukvUAkBN1Sd1+UKefqrXMHPVaGtGIraHqwuEu2T
NOefK1Fys23pN2DhkdRQaRj5DpZk4Ym9GPcPlvWS3cXZnU7YqND4VMijOULUfQlrV6SVxAbhKpCi
SrfdHJTOF5hRYkE5QYz+8NoAXiJZ/iZG2ZewFj6eLCSPZh7LcGI7RysIxJs7yaNyOwAQgoxUB2mF
3nW+sAnHTq05WKGGjBLR/gFqsM0P2Hm6GLRUxezwY5azuFXo0nE7EF7vwwDPTuOQ/pylRrkRQt/U
Wa8Uc71hnpUTvmikcrlsQHzRoqsspv2RX8swgJciwLCWiUhz1r5iyN4ufG9bcUl3b33l+mezKMSO
S/A54901O/IR3vj4anXAwFewPhI6gsynPW5nYPBIOQ9YwovmxURLyV7rh+Yor8Zh6Dr3TbXgLUxt
kwqF1lPUJh2zhP9aYK4EWfJ4pL8te6CeXdv1rIX38FW6FwtfRsTmlMkvEbCfb1V/YxRC1Q8VBYHX
ApFJu1eMbetKWmI4Jbi4SH5DLkCxUkmeeEXSh34OqiZl0uCjXSZJ7FIDu/pKLfByqsvXGq/BzUhU
ednxW53CmDOOtHzS+SyY80mfG9/G1s3+p2f1zpJTDXx64GszT5zy7a55+9D5k7JCCzw9g6TzBk1y
9O2Ktb10mPjDavty9laMflPBuEWtMGG31S5SVhv5Sowe0E/WoyJ+746bmWCkoWDDBE/z3RDkEmM4
x7WGTWgkQ5ZdGQf8h5lTuC+MRah6Q+OjEUsIVNdo0HWdYSCtggmuW+xttMi0JXtschPPeF+pj+cs
V7I5SGpNkt2y2I84tjhI4bUeDFhznQACiFFvGeJb13e8PKMYg9z69+gXddEkj2I4iYncrjxxs7M6
UkXKqJKNUf3PFGAFd2Jqg/Vp55kdw/ggQczZGPciLAsJotQMPb+OrMxOT/V8yoUcViXqXMTGYHVo
onSanX08DSXFS1UEnn2L+CfW1EHto7u4CqM0S8i/J/qHfptqz0rRjvvqxrPSdmOhTSmnUMM343yJ
7Opky4e1M0bYHdwq9idtPPrxk4MmqFECuBlh4MDMjwxoFMSUg8xEgjjMiWXPm2Z2yiX/Z+CrgvsG
7lUSjQ9cKJLCCTmq9PAJq3pu1No7M5LQsSBkCoxtoeh8S1Sryxvg7PViVxDEk8VVnFuoAxVjjB2P
xo0N05zJp6r4OaDLaEH/YuZyXzGXwN/+9AWFnMG2TSxr5UnNPdpfAWE9dnh5E7aUPKiUSIOZ11mL
QBW4gRHEO0+RDY+nIAzxb4igpmwDOzq4ZykL0qJUHp1kY4yd3YLCN1yIb2L2HVEcAmOllF8EgnXK
PRGDot2BTPUB7eb3LuR9YteqEyxu3BQwgExlIGfzJGkGwYlgkZtPb4zAecb3iI+fmk7NaSF2nn5/
0eH1WpHUd2Nu3EcZEfqCBYIJuIma2srTIxOTH7vYBB5ycSydlbd0KeycNAfVxkdXSqbOFZUJ7SMo
LudGqckvAXBT6aOAC6WDIxpcIgrjQL71fzJFxs/FpOb32pvc5QwNqP39jT7z6c7fXp1QlYUJV1R9
sg/8RoyRRJJVZm1K0F8Rx7652psYuXQS1VdaCdtDEV9DlLLYX+E0I8Hcs23QXpKqcvJVmtoNDpt0
lep/bLOOBdpfwtZBlODRfIrAu6+o3DXC8k2u06TNvOZTy8eUkf+rAPJzxxLMuQywJJ9aLglQ2rqj
YOGK8bUZrmodda/KYooYfVR60Ou5tlldei3pbN8UmrHWbHe46CdIeeX4IwjE6X/Oy7YL6rjP/2QE
WJpsAhV4+COHkZSsYyavsWAewJ5APs8x4yijMUKw9CiHiipKunRSsPTFpcWnLWNY2ETo/0PHYc9X
waQ3fDaCxQ5+EidtrFlZ9STlHZd8C1FTolHd8bR22u3QGXVdWpETAOGgHth9ztapOqNEXgPcSAb2
fLHu8bpKYzCLpUFP8x8bfxgfVEtCqm+OkS4Ph2vUqLJFGYCKC+KfcW0uRmq7lveqybe4NRfckNu/
MvB24tf7d/rmtbuw/hsB/o3lv0trMqDTQ/Q/SHaEwoah+twAnezJtxldD7LyyY3UF1J86ymS6Sk9
/vNBBAyPw5eJ/w6FA7l80pqoTGM2z0k1rCbWYJE5UtRz93O6IJKdNnnOvV2NPOqnZSyJP9MgUmPN
tvovgqSBUqa3QN5p3hkYCCt5siaJ31ik7fpOKbS5ww3HSgiV8kAs9UFcyh/IQjjadADtHQXkVgT0
6dhVScXQWW+qsqgR1g3RjzZ9pdf12HZtZdNhujmUsb4paYI3buw1fuTKQTDY3d6YpDLHuI0Bl2IZ
yqAMyn4p0eco2Ye7xbgntRd7rVMD4rGKu36PYjiUuBmbkYSTjirBb2koOKAaYgWjg3CZBWBSXfna
NT/BlncbN0Gt2EbYRW4wOYduSEq1O6UyeThxlgo1qgquWXn7b3c1Khpf7bnzDkezO8rKc4h7LQTS
xJOwNCyfZLT0HK20MsrHIrBfeVvRR6xhOJg9qUxdQzVIm03lyTgqJaDUxMEW52/2Y+ntQTU02WsW
+yyVDUuwNr1C2PlL7dTqN7IYLOcQKnMRc0+QOp6PNiJ63md17OEboD45QwhjX1VSwm4jhwWSKPHh
FgUnJC6MyFfG2tM6oXpyzOhB4RPMfHe+gCZU8179+lQUGogVAp5gsH5JC4kEzn4Qbrgtz/jkR5Jq
vEBoWDsRV954detbELblI3aXyaaTxhJN6y9wyPNW1+JXNAtxk9qY/nxcUCEOrFNnrPBGJBfLbU8J
C5T/ZVC5RSeAxB0kLfUDuCWCv5Lb7A5jJOJrjhpLN/OapSv//dJ2aaP9ATcjXrwLLscpR34yUv0v
hIUDbLA+gSkkrS4GbR0wcKxkSKY5hoevzvqptRDAqILmb/E9SWJAV32YVUC2FZQaF/jDQWGyiS6O
ATGKMhpg2tEjzs/77m6OGA3U9EO3BWcD/pGIYkxn1+EpsZcqJMKnVG6miVwx5wGcH7p8h5Y2x606
hyWmfPdK4k26xB0IUZ63yQuwnQWrfe+dWDOTRKvOyU5tpPLb+/rckxC1RvV7P/y677jxpHhh8Md2
rYzmlViFE1IBl1k6ISE7bCSdsIu3ZWGHi2ffTyCTVjUK/3uN+QlpaCIGeyO85xqCNzkzrafAOu7x
PpFWfzhK1UEm/MJXIX7L7e4J4QAy45fd3Ifi8avg46+uuIRQogTEwqKaA/s7YM0t/IxeJh+FuPY/
JY6rt9YS2nNUxlhG2ehXGCvumkbjvHZQWmxKYbg4Uv+vh5NGlW4X7s9vGvdahoUvXOj0WwQPqCII
Uh8Cv5hhmQvMw8m7pg42oFA72IujXSdPGi52A/veScF8E1q8e1t3SPC6gYY7wx+j9aJMDSd9g74q
N7neS60Q1WmBT1PiRnrjKVts0bu+507qy8DD0Vsfzu3KvGgU6iOxW2cpx+ybx9uPeu8hBPSJJecK
ie8bRuAOZmFjxc+4ivWzqKzZeE03LtzlZy4ArCAypqH6kaaRBVGrGw4bjvo8VL5iKMdcqGVrFtpv
GpWPvEr0XUZWZ+GFFaU2q1YSx8tCr1VuSk4WlKYqwuvzoOTUDWXnWo5ZRE/9AmVR0YnqzJ2dAoc9
rnmoAB/1nic55/7wdUwg+0Y3rMtySaeh1+7nsmyH8aSEOg0tDeRqDzhaTBDKfrDW/IOHqbJINWi+
9WiSxpIzoriKAstdADGF3DIJrO/6NKolerPyxLlJkYxOKz50p8KP1junqNREGPDo+RF4/AKa7vNT
a7iGkTRaFyvnUu1ATgXHpaSaN8Xg36uIwQTRBfaHY1sgs9ensX4HQwOV9fR72pAn0MRiS9CxHduF
oKaMFYoKu2g9AaA1oaR+ChmC753v32TpgptnnGgWpIdT5vqdvuPxXFqEIJfo/FjLbcRA60EgZ4/M
gMK/YfF7hPdZSF8cj1TxJWeQgzwTc2A/CzfT6Q1PBaeh4pTkPulbPm9AWv39w8TT0cE0dKa+4j/j
ZybhYah0oMJdUAz/12vWawf9gRAKHzTjBkS4iaaFli0Iv/MMhSev5nWBakgwISIpdnNs5pI2yx0j
vFGUgjXA8Vscxt9Jbfr1xyP/NLnSVz9mE/+YmVTdjUnNsEne4M5dnF2lEP5n5KfTGwgiSAcv7RQO
WZ8jibNyDyyd4GNmgNjd3j45dRXylad8Lh53wfLlGP7rd5OJ/x1KYsVvMLtBkkY6SjCdXdD0dq9U
yiffybgCkjYFJwxy+mfsBpoUJudHuFyOihPriOIu1neZ0s55dXpdsld/ZuuqqDLvnHiKe++ov2+X
wmfO9TlZWudUREL/JL9/fyWJDBazpkiEdS7GJ/sfcHKKg4iCBSkksZhKJ1bEE3adIZXokbSXg8Al
GxclT/MqDNGpBMOSbYGMELC4JZYQ5C1nzwR4rledMgIY5mTdZGvyj+lvbzrT+KyvGdhEiD+SzQoC
p+Qoof0PfsFe3cyCfT80QpQnmhW5uFzhehP06VnONL6VmBpdFdhl7OcdBWR72ma7x2NoCiocwNF0
uwUQ083Ncqk/qcv56Y4tsG0s/28uV3KOJboPuuowOhwQ9tW439HctL1J8ltLeVr/TUcW/riSze2Q
WcxLZM/qYUz+kaSucOEtUOqINaUVSj4QzK9qa8N+NIzZgaPT0vpHEkM0P4bCdFpKuCXr5iOsrmbL
jt13UxRlj2yAgyWJRuZKs85DAE8jA8IY/zERxM9yoz2zCVxpkmXUmYXAK3a44rnXPW5eqUqlHqgU
VOk36lles8gQeOBlHYGqoUJgf40l5G6y5ZlSlxsChu4bCMt5ZuxYZO2/7QpuWWK2chSsLqI9mG9W
35paDJcRD3b/gnyxISojPBegeVa/LrZS5IrkjfxXgBGYHcIWQ5NzjkD3a2i3CYLwajOI4icgxTK8
W9P+fmsycJkCEtK64Y4i9bpB+VkQa4hNFACkFe93RNe90ndicDLNIHZKOE6MC9xuxgJBByOLMKLa
TZWPbvSDOD3mM/L7khYK6/ZQckKgyz8WCU9baXTE0g2I0ylqfIhi6QqY5uU3WUCSTRFl1oXuzze+
ZmywwxGfnNsoTro0l3XICtgvkIBrix8v92GQLwobIFiR0SnZHj1+Ygp6lpmmRf58q6LzWogSy2CY
47OcaFdq9771cOyappKvpzTjnaS8k8VZpgVIcVF5JCkcwOJ8VWpfVKB4HRjbbb9UyWbZq9Ea/Sak
L1GoYAlKrXF3jy6sDd78dH7oELZg5gm3WQWeenkcueJ31eklvQ5IiWX9CZ+D3IYs8vbq1tw7LA71
ZcBLCVY6ZmLffHrdSSNp2wiRBJmyDf+tHACRvr7rb5LdGSiKgsmiJp75UC59S/a4vufXnl2x7Asy
hxr1rZ+8CyrMiL57TIHUsuKT+FeVOL3kzZpcXEAM9SV+yrCPDCZR3KhtAIR7An3Rbv7J5eFQH2ks
b0bOGjbTU+TFi568rjwaM5SVpLfHBj84Ev8EO8U2lFlVLTRLMspYNY/Uf3QOC2Iiu9JnHXYhVieA
eVFjiIwM8aF2A2G9ktpeuIlTBn0TmzS8OhUhyooIhY4ZAWhSKvL7iSR31K3E7bGla1tpsLTc6a+Q
8PsYdaK2UdBTF8fHEy2QTfXnoUJIczgDJP1Sct/VusdgQAXBxhFLdRzTQdW/4ZkAG4Uk/4mlHfEV
CNaP6FRKTL6GcjXWLlPBLa8vUF7MTfULzh1rEJ/cWQ2+8xIOOKCliK3BYPJrc3ZtQjhk2CReRCup
NJACWVTYnYjdXDYTgNMAqOgKICARrumZymovANJx3bwSdYNOyYtXOxprE65BoJOhb1ge1B2OQoAA
V/joYGqVUP8O3NXw5ba9Phr/BK3Lq40is3f0TlxRAKY1DZd3FL/wIHZtbPQnO8PnMlHLqHf/Bxet
o48falYCG+PPWDYvYbPawMQIQwyh6eCyJaaq017fl8/397wP1JM7ZzAEoUwgYrHUBMbduqUG2Vb9
PKjYGmESGIA/dQFIXpPlc+EU7eQtm5VzL/Gi4wMfHxaiuoi1DLHMwaSS5vazx02S3dl4s6tsUsZo
OufnMsLOoX1PqzPG80PaZ42re2aSURRREw+37+2UhMwk9taVsL/U5uFZU4gNJxP13an/aWqT2Yjn
AVAoTjifYND1IGKB7Ex7Hu8pjkpRbAlXpWTn1TUxA3HIEdFo3KNBRq7WkFexJqnBXr1FIS/BNYhF
JU5U5TLtiMA2VcWjVqf6Mdy684zgSBMq+QGySNGF2O5AlPM0A2dJwUaUczip9b6d4ECsuNKoLJU+
xYYARc+WB6f8k42hxxzMMFGu+Nt5k0z6yq6HhNyquM1X0TXhgSgKOzLDrEzcUnH0H6RHslDDr//T
qz02zv2GrJAbn2Z8p/MlBE5M6FCnXFHv22fHAhCPjLxaKEibvYwpD0LQnHllphDgEsTlH+inm+Gv
Vw+nIzmi7n/Za62b2G01y8T1EfEWVFPRwoYtfpiks+HuOdzvXXy8sXLXVifWhQANEFx3Cfal4eOg
8LZp4/ZpBF6oor0IesuYAtLC1ivXU4QmNRaPFvsqwBSbFSA0Pt9rXe+3iqEgxu0LbAD569A2awR2
ssWrUIuo+3OdzPdOWTWzO5+RrjYkRtqwaX+5/48VFy45fUOJbRrEv1gGjxJU8Cf5HcXWSXZRWIhn
Ny3Rf97fIqNq3uFFGutmbFqFQC7apxxMPpiYyLJMN9GYDXdH5dCJo/3MTceO4pqwc/u5rpEZ6CE5
tNXBhws5YWoOWfGOBinNsAibOwqKQ5oPwnDbRIjSxesbWoQ9bIDQDGp/2GUiLEalndUv9gwQiOR7
K2CmHkQMklO9VIZAQ06AzfsvdjCgmn1/QNkvPJXTazZuPHb3buCHlaYJTxp/eKueYbtFdM0SbXk6
Q98zRPDYt4GDuT1lyFvvCUQulftqIs1Gu2lBzjOdw7cXlenZzohi5/czM7tBdIWUIgJlUaoiHq6Q
oOhdGTfbto57sw1i3EpNutZIZBRdc2+H57Fu+Epb5nuLRfWHrdCZOkyk6K9X5r+RnHjnIkIwco4I
9/nqdgJlTmd6f7dO7OQmLL9qHNUSFtvNaI9gzQLQNZ33lmY+ns8w4S26I7oLu6Q+1xfD/s5IsrO3
aVVNtdl5IJ8n0KNc8HbiMiGV0+36ac6VsE0USoGoix9G+BEyKVxXquKYsbYqsLsCUvmxc0e4/UIg
ZPTGtDXgjI+48W2ZKFLKHTQVCgxhuj+9yLja+VARTTbdgySchT/bchrFMUMRiQhqnX+7iLncNsfE
cdZ7MQ1dBWJMIBd6fxQDw+mZek0fPIYns/baPZhIkrE98aRJhkKhxTMdSwlKJbqqGxw2JRsA2WXt
LkblJwe9QnoXYC/A9Upitvxl0nOCVlHYigkL/qVPcItyQcc6YTAKXHDaY4zjZFgKP9TxgwC6tpRN
xJ6UPilD3D8iL8cQHAGxv294WzM/PvrKsABfNWU8hemrA/iIbf/kFn0nHIAv9J3ZxrBNyyDkMRAA
D0Pv/HZLMYZ97go5yxzCb6mZosi8HM6PxY6lV0ZnePYIKGQzNBx2egJUiXLIRWzCyQqMFBFZXhXv
SY20MVGNwa3oFeDkFHaA1tzWYcE4FX1dXHrfbiGL9sfzcRI5CpQFl9T6jZdw1HAVuO9lB1uWksKP
8G+YPvrnkhX71qn4j/Pu0aJweH1LbXAgYJmb/n4OJiHrcDsE9GlDqtAHbQeMObFiVe4+DW3lVWiV
4jivZnvc2WCD2rb4LgQLw3Qc+5YTBbivDhSAYXR43qaRsqjoxUxR43O71j8QDec2AmZhwdpziFIH
hQx95eCRsu+wM5ElQPuiahQIcOJ8J3t4Y6G7n7b2XzgvNvobPbARHK6Vy38SzxFRh9btzN3yEG4D
OsRr5AdtQFyT+njPplREczOCtnZrJeHDM243p88eKl5tmsSFJO7WkqryhH4W89Awj34VAmzGEh8q
H2m6mk1rSwq/EI0ABli9M1KmE7n5PJRKcWqD0aqbaw5qKnSpvAt58dGz2D7R7O8limdJlNuwo+i5
7HYI3hLSA73LTp9gbzeKC3/suxSS8FPpRC5yYcWoA98WIoOCZ0GQWVGLBzeokZRMC9nBnA0zgbnl
QHYEuDzdsmW32JEsRv9+knkOeO0fjMvYzBeVsSKbyiWWOW9T6FCrqXd4lk8AKyrTDHtzCHsPpCrm
jTZgNMiAt+R8Z/TR6h0xLrn4uE+00V/kep0tbVZHKaejpstDC6a7UrTSSmKWgsjPjkbs3myzq0UO
MhBTqi/0lgu3vtaxWhR/pwf2aRHUs8ToTfcfn2Fst0VT7gfZQsG6KK9vqzgLJnVKjiwUHX9NM+D7
cY5DNWtdvvGT22xC2OxY5hpLh6CrTbnK8HtI+bmJBnGl9cAxKgzl6vg3BOjESon9dNWe23b/ruY7
yVzjS8qtHycuQCtJS0/cujSJ+e60GwcRGQH+r/9LTcgb4ag/XsWsmLY0dw05DTWIsjjRUZ23iOxI
8hEANPwykK4UUmO5mwilfScuwsZiSYa0rm3mmguOn0mAiAZK2+meue1TyQQIefHNiMMl8qagUia2
esjlasq7WPjRpayAT4Io4s0BayTXH7ZDKBWEg6UtexINWfPBnAbCOMLWHELgRFa4t0WZ4ystd2x0
eqqFAtG01wDZOyH7bx/POJbSoSmqiXuf20bTinKCAV05QGv0gqN89kY5gak3ztaeLStpcjV1qYu5
BVVgjlx6chweipJ8DV7ZPUgeRNxOv0q5kSuzORMU2RLD6vbvjwzp7j9MZTl4qfKBc6l5+KtYb72P
eJZtj8TNqmMf59m4KivXLo6QGK+M8wArBCGCHeqR+ChM+X3TRe2gsZQCy5HL8gOxfQRmWocjT/Ts
5/72Ee7irx80Pq9he0YqmQxquPXxPqfMARRLSnWI79LpOTcxodIsZ0h43ktAifVybl/RRV4/msQx
geiLBtU6/yPpqSrsYY601EW962DSN8K6wiz1GAeQ18zV/hrT1Eit/Pur4teSfGKUzBtfqOzVVDvD
ymGM43rHd6jXGUEKJKC7qDxicnQVnzMOKf9DG86HaKHHiUeOy9H4IgjGBWgjud+6P5R3QM70eh0P
KvT+jqfGS8YZZPuvEvkEuuDL9ksyiI2McuA+iwU0bx1wqINJt0vDA6olXjMLP5mqLkTlWa/RnqW3
3O9ML2fuzVUH8fHiAuhIkpDeif74yLCmDtKTW1sZ/3ju9jp7zDOncl20qDHSSmDkAuwd1OZ3COF8
4rpIvKGAu93e7braoXE2Ml+p/bba53/d7b3K1esfZ9/wJdfPZPDV8Z0pdlK09zNs4sK2EpIAyQ6y
yc//7hW0SctAdI9uHDe2TtFbZnHwUStB6M9y5rryvs9/TmaQdWPuyhc5Nt//iO29MdB0Jk93SF9h
Ad0laKUyH2t6zXwZVOOOr9Ubv9Y+u/aJRoFSnX3XfE//z3vhnLO7zZPRAFQ8GYF0jMAhCHKsvI2G
+iNQ0IW27mSy0ocTfeOqF1TWY7+VCtuZRJbN6s+xtg68sLMavJ0nip/eI2Yp51IR6tXEv2qnV9WW
CrvdZeC9Ip1XWslXyEtbF10z8pt7H/UgvIXSBkTmfL6B+2tz12Bezc8wJ0Zo14FGB4hD2frhWZA5
rTtfDOmUhlmrCd2H8QOKbTkb3TxxhrXxO/ECZ3N1aTr5LrWAzpkCJoOXFR6iLZ/H762mrrpsCoSP
MqzgByLrhDwEr6cQg9Ba+7ExP9JD4ZR/ECklFqk2CeqsAMWH8HtWiAXzBhCAmYV7np4FGRIZ3Sh5
mB1pZrdlUQxPMdmofoTemB8LdZeF7Ycd+dhiEcpFxcVlwU8ap1BJfQwdqRA25uo4VSzxRdFCEZbf
+aUURtvzD1AB0mUv86imS2ASkXZsLLHZonAQOqINqL2ywjtwnzO/GJZyGVfhWV7NyGPVCi01u5b0
QKq2geWOdipeyASQg2n66LDTim3Aq4tpn6PTb8hnFhjBr7etMG02dAkiF/kd8rNkFntE6XGqMudX
YdGkbzLixwjL0LDDCFBdLInUrFw1fdK4e2lFBeRP8GyG/vSCY+Mk4nz6UODqBubn5W+aIPIGnOWl
8ix/cTOBMsocnlOw64dHlB8hlUJr5/FpWXyunwEa3tdeVSdNe9OCoIFg/W/4D0siJtbfZJnpLxeb
+3Caz+bVl/IoLEhXguaco2JG7jyEDE4jmjT8JnBKX1ZJs9QjKhdgGFLQN4C7nYcul6eM3HXbcs2K
YxSd+8UCusnTQN5vj9JXPPMlZCnZJ0JLTyA5DlAe3I0c0wBVHhmLI0CbjNoOpOG4+hqThEvzhmZA
hDxZ0hxnsZEyERK5s00i//be/j3hy5iKNDLRTxK0rPYP937wsE3ZqY8XmJ94ucdCPZOXBheLCZHz
bwgyd+8vsO5yFQ2TQIeXBCZkqZrCAXd2OBJ5+N0IAA64c/MtDlhCwj0j3Ffn8rOak5lI59Ce/b3m
UKtQJ1008DI3I+bWrl0RkuabTpBbU6JqXMlUXiga38SUIuskK4ZiAjVMcddHEll4y17OQQO5QikE
7eguF2ldkqKtD3RHy0/iQ4pHX717BveFZkBVXn4OxDYoAN8sWb5wGqOx0eyS5pciIhInFsL41ES4
Y14CMURBZdm8Zbk8GLNWzNBdY48d7b6xWNSsSANpqbelfLNO7no4/+zqAUKFC0vdmfNxF50w+l2s
NJja5nLr5ywK6nRiCky+2HVT+MrIIou9ghpvNQSbZigeiN+nOlDgRCbCfT5q2HGlHNKpAhcHBhrh
/h4b/1+A5VKEWPjGO9+YOTWrfcrXOyV1a2PMBUC1oy3JamHkHUOFTu7sLa0scn+IRUssT/D3PuUq
zjmTHudHjBFkboBNt6opEJGYEiRUBEDyEFdYFxeJ+S97hXw+Fj8t/e4u70xB56aW7vOjhvNBp7lc
eRgNxSGt+A6X3iiH4I3VZ4ExjvtCrXUZ+B9yrxzSVuFL75VyCgnb8o2rUAyjz+IZ7FfvrJ2rz+Qo
umv8qaLiPLDfRDWVa2NnOYNSC7Y+Gl1Rg08afw9HOi4evX7oYZa/74+33jQXCtk2Gin2H2ZLBIZ4
0k3b66FEZr+WpHrwf0toQ6B6/8H6PSYsX43SG7I7CqtlPAjej5/dCsmL+WC+iErlDGJPecbNITKp
QLW/XocaY2MgqIC4HbC6cxKpZsWhM2sVB8YarOcV7Cm6JWTLmFsOl4rB3lC+zGilM/fLoRnaS5Mr
RMMvk8UPKrAyBrT8zebQPPQEJj3DmSFNaShKAH2p6flCPZHDKwoyGX9ehs6wGJM7+Enil09GEL+6
l/nRGcOsZGqwd8ARPZynwAZUtAHhNoTeunW8DvOMlI24WjBvwtEsLnTwUAGwV8lD/AcTKpnlCGuz
omhJcvXY3gjJGGKFfOw3BdFDeMSWgEYelSmrcKruIOm7iuqY+ruc9xIKjG+ibqLeNuLziR4luTzy
KhKFrmQh1rPjafjpYLV7eDlVYDxIYULyb3tsierTvm2Y5LlV+qfkzfCKTu+Zdm6sF0e2kEwPJd6+
d6lpSK3LuHxN3UkWf4Vu1ti94Fc7vtZl9KuejomejEt8nn7Bu+37PsPUrrUACUWD7BWX0aKBPKcl
2wZlO4O1mFqpgMx6JxsH113432MQdJaeh5mKMhNR3fBpIJXd96u5INHJtntrH9q8MI42TJ76CCWJ
n1UkgiAfKadj+CDoHei5S8io+zANOoziJgawsgMRsZE1lasE+g9q0zuoanY4FoCpBi57qscJOr4C
7RDdCte0neS4S+ffTR3W6rFeVzV9loACIXcGimVN8/0ehxpe7Y3DZV6csA+0hjSlsz8q38Lzci/0
/PTuPWQaw8AJOF5srWuzjVd7Oc43dw0af76cMdB2jMt8Sk4r96q88Vo456g3jmnQPRUureZAESY4
eBlnlbgP6lqaHGLQ0sBtgx3Xbt58OJuCVhYnEhcFxTqx2ESj0KorRYhLi2LYs5wLZkayGSBdKBzI
dXO7d/nFMtauTdboeOL2vtZFXyC78nsVaI5i28n0SOWHrlAcb+28dITjeOMEAq4q10dU0kaA1zlD
420ClHDdrwKP2mlPIfIChzMXW9ZC034spMqnK3UNezvqh0Z92lL1xmQ6HDMYRd9G2SH7BxDUmTZO
WlirAj3I3dXDhWtZ2nkaYMO9hyoJ+bqpV/yEcLD1eRFMyY1PVSb7V0TlFdJNB8xVhMVCT+k1KcOJ
K7DSl2dVPja8lEvJzuvIF9jA81VGqZmYgHpbwJ7rWSbAaS/w6DkL8ZV685khG9KU7aRG5tUkXYAv
GQ2QvEwwW0ovwQffiE2OH3P3kXMApzBvIbilLs+ndJqJLsYx9gC3TqTj8FwFjV0RuSsqhoZmORFA
Hbqs2xNf3GZvLuZ3n8f+qpHUlHToxJG8dqb5RVv136PCdad+4DRh5+cMUO69JGx94Q2iw58Hpogz
1XsQoC/kptEtB/wjS7DdqNzkz7JiKDFeeQBlZvxheOChPjhuiVBLxcJQGD/s5ABHv1urOzlPUgUv
22td2jBGL/xa0oL9C5UaE3I6jQ5NyZwLtwFSWiApKrowJbaBb188lE+ahW0iPS0mFr4cDe9/n9Xr
zO0LOnhcLn18WAhWRrUIMnLO6I3sH58hLgOmmx4amimQzQ+f9XXq2E4X3JPTrj5HfU7eEJb4ERIu
FWKEKNwLhj0w+ud9bPGF8ee8/r370u49xpJwTNMEc3Xsc6x6rp5zbWkEnvhQHaTqpBV/wZPR9OZY
2QHyCDOmusxw2zqGjz0Xqpv+hqLHD0qK1T0J2g4Qh2p8rAKwZf5x+485GCrsvBXGvc8mRXQ/GgmD
aZcGCxl9gjjbdL26TUFzFgvn1TbCFWyjLX3Dc6YoGoXKtFP2Z1+57EcfICwpwqklELI2brGpMxLR
bwYWFd6BgYo/DdxHCA10cydncPQ652tN7Mkbjgivg+x1RR/5vhYgJPH6ajvAGjhdb2CjNZSRKL4o
wkMggrQWrpVXGkdk6wjPCRUBGKk248s8G9lTlhvDbsycSvPLw6uYMLkvFiWuceagPj+0T+NMioVR
+079a+n7fCgPDEqig7/1b6pA/O9aeJJF1ip5amnEaWGeIAVQoExBzi/471dYxJCD8K0e6J8bZHJw
ytpQprejz480ZQpzAlyoMTWUORQ+zC/EPjZFGabZ0mNlh6TUQ8InRXuZNxLT4X3tERN3yNcgwiqa
GAyawutaBL9cptuVhetZ1qr/WFaKSkaFs8pKHnzSULII52veddJ5lYu/cq76X4iZMAzQ8BDwXTlI
hVdtoVvryH2Butx2GhMm5R7ZVzwuYVvauM0gqXH5dt8LvxhHvO1EtiE2Gb6u40vF+xgYzYX6EzuY
ndlUzxWWQT2zslwlGuVOEetA/EQgGqMoQwgkd7qSqZbuUcFZAhWFuDVcYT7IdKBOH3QH0X063Ixl
eo+I9h1jGfXzfNRzlLx4I46s9yXiKAPFnlz1/KvYz445x5KaFWmbQRxPWd2w135F6ft/sQIfov/W
aEqXt1KhoUmlJ7vX9mWrQyHdXDeSZO6ZjtXQg9wRwx+pCOz293mUCqNJG0Zi9mFmqBzF+/nd3/ku
AERWce68IwVJM3N30Ji97n9Y5BwSZVAOYp3tFIZc9+NkVKh/JFTEc599LY4v5VOJovHfrXji9Ghs
3qI9xCsbnUsu16Mnt0l6nTKQfdPZWPUvkKdmeKN5aVdkcyIrEWZrpzM5bksIWjT25zLE84iAab60
TFYHADCGFbJ2+hx5asQ9qedH4qYsKXcywUytU/sw6GBorkloHMs7yASaayJb0hQWaGQkrl5GBHpo
5SOfBgnqvxk7CKsJF7pTbArh6cbeTkFOqqIjRMcabf70wRw2hAHFITtUulUMg8ZTnj6B/D2SSctN
wLWBIAcrww08I3pY5LW32spXQRHDSd1hQXvpSBZwCNYx8XrKOV7TSbj7SNSeCuzbxm+88O6DIsFH
J1l+mJn6yCvWfXGE0dLPbEFgq7zXoMzULMkHrX640PBYcuoyY/6+WHnoYxxsbYkNnZLu7iSfLM1B
QudaY4RUGJklCe+9KiTnjTucTK7JVCblGxROIbyo8WA5PGjM+9dbCTSwy+tPORJr90xn3GnqQ+3c
dSnRqz35epUqiIf0808As80jXYFiWUWIbNNvVCHCYUqHNlpm3DTd4OtByfrsK3VHfRev2A==
`pragma protect end_protected
