// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
w/EVVDu/5yYqiXbuOfe5gibVHwFzIpSc0zBYk5lkEUXTTJEaup84pJaYbVl6UeNLU9bxL0G3n1nR
hpxvZZ3a3u26lNLQY8Y13eh1MzDOWKWdIv9SVfubwAR/L2Ttd5ebSsGQeVmc8qb5phaffpeVUOsU
Q3BoEmA25hDYgN8bMlCUU5KZo7VHV3fNQtoyay7hPoVfmwoCrPabbvivIkJDx9/dTaUkdDlLDIxq
3YpBD4KsoPwFy2bx6JSnj82T27VMmynPDNR3c8x8SQOo8oag4G0La3/21v1HNL73vpeasmagXSdo
E2oc6vFcr6syqsFWZkMeZX9P3IMqjb0CAd/56Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14016)
m2wgVrhybmU/vnqgklHSnx8TpUBebKiQBsDypS8bIXSZgzH6qDmpn1wP9+rgqZAp2HntmMrWYKsb
ML4gMmUnz/UZ1y3wvaA38G36GdmjXDdxWR7+yPwcZv/0ohu+GM5sVikV/wtMXOSpBAY+Dzo7cUK9
/DrvB1wo5Cpt+3tCM9xRaSExISe1r6qyjbLFmme6y1lxgTMHmMdvCfKERLIR1IqLHmXl+9alPTwZ
gT7+GL5UVBxxXZAUg0slApNv8LAA+TQsBK6bjrrvbEVeU8k1fwDgzoKM9YMNCRV8rXdQliZOkOoJ
4K1MOYkY2eWDjW5KLzGBVmUTJYBjDOIm/n5gMjq0/BIDUCiqdRvINj+tSYYaHYgq3rqmhKNhd1RL
apLMn53XC3i6ELhetRCSEsN/ipiRR0VfZrbYuecugMMOAZAiHwFhG5/X8Ez4ka2QMgoz3WVMgkNY
VStUCj9OG2N7Lq/WLlmSFcbP32dXu7ojoFcLUzn66UCRyeyyNffYiuMV9k2cd0HWk/aMrx2iLAtg
qPOtoGdtxkiS1GXTfIsoV3AN+JsvopTfIQw82tN9Kx8D4lxwFjHcvZ9wUJcelW27+uLqcO006ngE
nLwCQdrhhMTIDJDyTMuZGk7etMOu/aEgTiG/qOy7FryACFFfUS1kW+Z7Rz5my4tawgibs+W7zF34
8SLx6mVeQ9VfeUBq9gObWhKLHQpzRd025Ux4PhjquP9p6YdUZCMxLDNIss8klnoZmPGK6ro/8hYG
9ascI33CgFV3yUEGG4LELafcQ81y1nm0pxCNV83HEr5JJVgOp4UO57fMk9ou7FiLe9yu4agZvVVD
BKF57eYWrwjVzq023BOkXZ4MegiUygYAAwB1jq4ZIKjTHOjA8loiH0cdXZDK+NprWMZGLea4rWji
B8vdbJP3zkzVL9+rGcQ2hMqCtbZlLGmJzNSDiPsAldzMIAoMzcCpRbtER55ikCuTta68bWeOW9rE
bEOG8f5QELcQD9wA7L23usd+kFG8SXJ/SVztL+WgqwObBwmyrVPIr5QSRn1jmUL5ELTD084veDC7
ux6De6FpEr0SHZRBvSW73FIy+e5R9F82OYEeBG0Wn2BS14h+VMLzG1Xu8U+PC9NjSiWsk/KBMazG
pXTqJm+0VTJMv96KrJSYCOHKLYrowgAxLKOG8cUkzxgYvOZwWfkqSN7tZtEsDCYiyrXkkMpZbH82
ZHj7hPytlJCBAzFEZDj2e+x+CRcYe8YLCMqB31VVAOSMcJMhhVHUNzC25OYmXoUZk2PMsXxnHM86
CUsI+aRi+jQrXUh3iOsFSDMVgFzhRndOYUdNfLSbe5SJbT9rJ+nFSCGz4bmf9okVnOnKA39LYGeU
hXnsKU4zIckCwjA2nWQpYDchFVmKT1o0jhgQq/GGWG+ZfWOPqKEjBnPNvrXxdAXjJJdciUjowRR/
I7Di2RdiCbKncX2KKxpEV9OEVJlXZrU97lp83cPrPpzRj02qXCqwtEAppRxa8L5ZHsqUS7bbFHwg
kFYiJeJVHM97FGEcj/q26iEY41hffsQDIulyHNUmLfR4zxhspaW3hNeXqQu7eaD60hTdcfrSATyv
pI3xVZy9HPjM8jL7BKUxMt09jIxFI13vMKxAIyVMdCoOBXl0rMz9YJJe0dte2wZ2/vhYJuW6Yh5x
aOuo6nKm9QhI92JCQ3lxuOkJKdkVXbaAEnLcw9vdKV0BeyBLjnK35qsSt7rxTi2TR6KFDGXDnSvj
KynnxCinHuBPHHOL5ZAiK1XH9MsFNKa2XYEwjElkluFkxIDpYze2g+ZiV8zxfZT5IIouCiB9urEQ
M8iCzvsVNm/J49sV2F2qPNEtWM9wN8Rikfjy98RUXWO1KFHPCAJSVyMe/wWt/YzG3K+JoerQcyeF
mm+UYJfaaB/OntSG7oUD9JLJJrh1FmAKlam45uncgv+mIVQx8GpdsbKEme0lkDIpBGfE+eFgeFPa
zAiZ2R5zq1CFGrZjk2popQ0QwxMnqxVldRUZw2F0MyD0tbyF7TJPyXGuT7p+tRRun2Zc5DupKv+O
FwBh9V97+DiwYK/cMCXftNsOXq2fqB+PRXgfEoMfvGTpAI/BOuwylws6FZY/8rmg4KFLF+0dVsPo
IM9mEKw2is57JVR3VSVXENL4xt5qztDAGKlSoQZeu9hAd8FFiA6FihHB/tGLPqT3rTg0a3QdaOmx
o3WUT2O6ue2F9sPXNcdSfIM0PUaDKC+8Sb+5PbWRnqn5ZIFPqTwfVoS6P28zr5mZousCXS51Fhjd
AUR/bHJUHTD25m21OTMWljjsxtR5XGDde4+qBU0MznhVwYpySAYvKr8yFY7QpwqyyktPg1pbBljN
Dcjv4TymLq4MQG6l889DX2LxtG2dFGAOPxOr5b2Y1dl7AVgLDkUu1ZfbZAmZ3tfqqvoxzhQBaIDG
opl0VHU+sFWKtuSsQdrI2zEvMVYqysJK6HIHA4TJe/02KYmtcdKIT1jTtm8Zg49cHZoyaaF300Sx
DgASJ8sMzsfD2a52NCYl3eGlK2Kv2InXxj0cKfu4K939R56tKxDAUygeyBMoH/4HSmK9ekg5FmlB
Jrq5RRBMu5rdKFj8HMVTtMESvz9+jp2PVaPTx1nKax+No9HQizI+jEmEeo47rGaSy3aT/dQonTQu
sqLHIKf3HrlsCixHlYjNiwvJGMU0EX1m1/MWcnKJFFJQ+0J0Yagb5/vORYJTGowTLGKu2E11HNGa
XwyBZgpZ9N3uuOtbjsddR32Ju6EnOAL3cV2dxKLTmwAe4mNL3TbgVHD6jvZErdDj7YQ/4P+Tp3Rt
lCJfE+2K+0vugtvtd4XQRjY0Fh6YxQlyoObbSh+ZclPvn8RBUF8JIEZ6l9xrMwOD6e7Pikdr7iO7
KYiQ1ERfKap3jC7p2hjYzzo9Nj9lia5a/RawuiM+URVmdhzzdiL7utPduBY0tKcqre5j8ZuVKLRD
vi9Y2LouIeUa4cWVcOm3IdFVcELSfEd1IDdxv8v2y05CJ2m1e2tlnNOEvEviA//0iVUA6+4nGORF
JZ6VPwlOeJ0mjsm3vY5AcYDEnpSnpRNbvIb8pVFa9sbC1ZotuFtHTrbGeIt2VzKeT+/F+6gz7tcO
iJBiVka2RKDYyG4GBlZFJEghgc0bBukbNzfFTV6uFERK5Jtlib+3KCZUYT+TkoJE5x6JOf/3MPsZ
NbWP3aTF+ObztGAi7JfwJyFvV6tfpiKOeuyoDbZd+wNrOTWNyfvAk10AiR6rbwLcmX9yAILcfjut
DugJ9M/I78B8GOX/lxoHeIzws+qzYI/lHT6WgK/+JCpoiP2+IaHJvuH7OL0A1+LZSxCEnslGV10P
jbOb20ArR+E+lxhMoT8uMNPQb/1/BG08J8FA5OJkcbJB2RL++Z0t5h39NU1rV+da+5UsOfNM5Ug9
FOtw3PAypNoSqa42j/jG1PMMyQuz6xBHTtvHGmJvM6E4kkd6Ntz4NoHbapkfZX+cBAK7rbfh5rSj
3Np77VDuZwFagjtleJsb4dnd4P0Nb7Bsi49Z8BeQt/cva7wnVSIqPWhpgtekTlqVvG1jxDkuVcnc
pUisXk9XC/wueIUHISHByb/dm1M7S5doZLbh4hLUIVqiI2hSYpv0SEXWVLdpgEu5XQTq7wJfbtPa
mM7GyukJfFiLmwDy1Ks6SlroMx8THh6rQpiL/dDBRgiEm+8gd67w/nlSzQqoRVPa+n0E/U6M3Gh2
SKcN4FfG5Jw7mbIxVEzkXVHdrjq5P+8jEg+sCyhjfEiJRnkOPozUvxNiz81sZtiqkJxYZ85FUFpb
3r9MF1JdwhB4p4ikAJSKWQRN+hpcQoqcVbADKXBgiufOki2rF6zM5tWKKzO7xW4EdvBtEywu2lnm
nbDL6tNG6LRat+MRRNd6vZGnmYCNJGvDioAm2QjjNSIxi/dZJ9HgsiGQdObbBgE0ICA8OnHvKZYT
qDQ/1RuHtyH5Dt+arxY1jF1+Hc0FCWPM2dOvZTokT+Y1qNGCU3fl8EO2CbsVJbkW1woE2XtSEsKD
Xzay4dv14IUi4QpW/EhCa/PX8EkcCrOMMFs4RiBxZNipG40AihMS9N6YhVaY9hdXmd5JiKVq9GgB
RUmppoW6Af7YEqpDS6hDP8PAZOdTHLGM/oLsEz7f/sGwLM5kQ8n+xBpOT3/N6FoGnleFx2fYWuYX
AftwNV9lJML4NnsvjLCJXiEwR+vrU5avZFLPkDi++SMATWaTvNwVeO6UFrRshSf4VO4IXouKgJPR
3rffxL/U4Mmc2x5UzD4ysmfa0fZUUgpXzkuPp2dKEq9Yfik2UHnz5LVoO3t32dKsfCw9YQo1r0gD
yRY2nfgbsf/jm3NiVSvtDFR2geVNxPEJllu3MDUAxDSrbDV0J0zzUERGloPwGX3fFp2gjd6TtF5x
1ATaBRixfbrYNfQm410ZHLS5bg6IuOMLfLJouCwxbUK4EiCrRmu+dTiQj3067W5Lqpi00I1MROaZ
6VDGJlCo8NVvWV9a0MlmONbpibiytLAKp9zi6c5Sg0OUj9Hh8Pu7gHFNVtWNAcUWmi5CJ1kYnoGz
DhSGMg66hnNGaJmEeZdmyDZnNyYhISdO1Dl7B/8MhWV2/Js2GBHmSaOtsUzLZ0D4Wx8KtaHquWO7
LEP/EAHfoU6ZVXgyLgXL5PvsBN/Z8FACeM7c877x5H8aZ7VXNh9dPVWzoRLa6MA5WRQebTKp7Z/L
9o0TW3H1MV6BEygdEQqeskjKGhilvN5K+CUJ7nq9umiEb+Vl8baMNEfrc4iHIbXWqePQxKHyr96Q
bRJPq7PpVGf0v5IE0xdnojnLzA46YhJfXzrpheB3Y6IDWX+XzemHCVpEXQSYo5foJMtJZz2Tc3/l
KQIZy64IVWCsf80E3memkTZi58E2WapTbDslhNxvDiQNcAgwiFTeWIqUwCX7E1PK6Rzs1f0tjE0D
gTzk3VgnC75sXejFvSA0kA3XEBMkRgElBSkcbrk+Fohovpcdxb0eWQJiOHd55wxFbsQxNULOtS4s
AhMqJJPbBCy3mBX4vsBaWfzIF2ZyeaD+2q9NzFnTwqHCoH3IYedtEy2dnYh2Al641/ZMsRm924xg
WuNfQoSSsgy0GBLTh0lH1g2iN2AH2FSWsc1IPxYHdkkt+ReAvIYPR80zTGojAZ9XWmeb9hswK7TX
8gMN/lq6kKPveMbKc5hkZzMu+FeFeAhpBaJaCGJjk446kVAcln/a9WqsMIrki2YYTdWnGAmPGlT1
H+/C7KeqHSygEfUr4aqYQ81gmeBEGqTMcRDxKkigBEQXdEh8WBDmz6nQJwagqACWce8HDnb9J66i
Fy3GjMjvlLP7fbVyt/aRrKIl1enrZNFmb4htHT6ooDN3zt4oPNADRBHcb1o5uMdRhyW2lCXZjGdW
gOMFtsswgvAdru1FpyNDSFH60JswYsj4kty7lMTViDFxifnT5CIOcb8vUL+G1z8eQADGhYdX8dHp
uuvQ806zfBLIUK0+nlxfQQv3cdrj5uiARuLgE7L89RiJ7s02adCi/TynwzqfhZWnqE8TpExqpE2A
tFWiVM0DIoX50yAO0Y9pjspTdbu5h0lZo4aH4R0jIe/ZLIbFeg+03pIOkb1lBcHGwyvtbMpOCCNR
3jCO1cu2633FsWbi1OoBvtgrJjPuchOHJ3l5CPX9P9n1Z87wa33JteDWg7xtuADDBR16nGYxzd6a
1Pg9V6qgSU81hqPxOt9Td+Zx9EykEBzw09HwjX+gipT4tP7tdjKJfYaWnD4kOMoL6lKvbLXigajo
s26+yIy69fjOLacNL064TpLhtjJqpH6uj+1f0JUGNtKFXmRXMep3j7AjpqGhiVX+gk/HAFu3zngJ
y0tISycR+qQNEMNuXwEcKapL+xfmJq8xXwWhhQHIAWQMEBlvsjUad3PCOJ39tuDgrH+KpJKpJ9Ne
nANGskeP+gq5lEAZFEPpG7QFiPjVl9lhwMqTW+lhYQNg1RvItMGjsM+hIhK9eGYQ78A1hOxcc9mO
TZ7SeRGuBY/o/Y6V3lyBb83+zNDzMLKlx1pUd8zhHLeNxKsbGpNRPgNPVt6IJbLrBEGaLkhDykxv
uikJ6Cl/S4qAes5YUM11q6wJawBYYxJEIOZSkKX8VnL/mDWUVNz/+0uO1E5fp3QlN7256lJRYWTx
5Av3N/G2696LmmR6Cidll2vMcgwPIu8TYlc/2b3wzcwXnQer0gYCrxfGc3x3QkLfOGZno2Y3nsXQ
xuX14s6/IAojY0+o51VwtoEnenmnHtlYrdLDoxfbrQT3vAhl8CeBV6OPE46bjPegAPpstY8KRN6M
dZwyC9vLzWj0gEM3loyC9ykah2X+pIKjZ75zMYaODOfUye95DBx7+2HN3Xi3NBn9vRxh0EGsU5CL
DKiKuwkE0Gb9Hhbx3t/D9p/txFw1cOVhCmJD2ZAtDBtkM52IO8NLzGsCN1nCt4zwIP59xODjE4N3
GP9U5MCP9SfGCERfVZHSznrEjDeVnbCsUQeZZYZfn166JCqQ6kiQ9cIUy8xbTxuwQ9tTKnitHgqD
qe54gtoYqbEbb4oI8o+VOMo3UW094+Uu0b1VbzSzIt0Ye7++Ybbsc3I1In0GtkoTJohNB9ULLlqe
lIKBUDKVIiFD9BOAb1MlKRxiCLSRx+Tn5499c7TeAvuae9yy58gCgepv7X8Vg/DHX5L1nua3Tu50
khnWwTW5vlHZJuqEpoq8RhJqxuxdpUU0W9EstezT9tnFKyJ5Si9OC5gM0gsqMReLbhJ2oCLGkINE
Rd7YSkxhZ6n/DleoN1vFzSsRggU2eEfTemMV8mswVf2NY5TZ6KWl4rqzSJ3SqTh3X66WGSm28ogn
6hUDr22dsTZg4N5AM9aRLhk3rJBrCT+2CBErcAYG4nPhhmg2TX4HpKmnsykP+1gVwffB9k1v5zE3
idZU0o60bAFa+0/zNlQrXQbV6bLxn/GCZarKGL5QLHA/661isS9Pa51X90ThUvy7VsRfEw4CQJyX
bY3ivm/Aaw+tomQqyZ+YnCiZR7vu4y3DswEFK4pfRNBkT+PD+BY/gXLo8FNR4Il+qSHHu9X+L66m
CXidqZ0KGS7WVV4m2tX8UQWczA3BRffbJ5yMEUWQIDriFyQRa2pEwj1wdT8ppG6pceOeqWM5Q6Me
Jgertad+gk3NcJ/GCRRT3CgHALP8h6BXGHe1YVW9VvslqBAj0HGq9eSXwocjsvpORORfqXBEMW0g
FXvU256wJJh2p0TdaMuxXoVXk3iQTQVkfRpqLzlIQhTXm0e0IuY+Yj3IaYn8LAfz1WE2zuybQsGz
0No3yBPvBHxRKwePQb5+9x/CzOmnRdwZJOlqf9IWpR9EU3yLqO8Vjj3y62O1dHSpmJ13/TXSfd/+
7PVtF88WinUnz67NaC7TpJS9H4j2CFPXY7q+UjODwJ0KJh/NYOBUpdRpf1/uJG/4HqEoR+WeXbPI
+GLftAyIDKea9c96+VOnbJJOlRD9Sdxz0q1u/YtktxmCs1evB9PT+pq1tpZKPBY1nvXQCOWMEuiR
xWE0IBWLLX+YGcAmia0wgh0E9y6aOM40NHrpGLoT2iIonZ6Ha+5jW0KB+IkUzexhd+rMm4ebJxPm
uAIh/2KQvKYqLsQKQDXQStvpjHiNi6Qx0B8DWV2kBZKe8lxoRjfa7bOu1VPmCfwFA/hoOdvUtzvJ
r6MTCBfTCkR9LmOUvhz8DOM5XX+XYUvTKvsCuZVQ5UTUW1p62hn6JjJ6szVBV+on4a1BnoWKlHzd
yvxowYfWY24go2PgCprkTw97u8QrWFnt5Z7JPAne9IOLsEbjJbRg1bznTomVgFOomWnG9UeXZLut
QEqmjcfQ9QgNF5UJQ2HOSAo80fDfdq47vd9ilgyCspENran8p1wN9y7c8KgkCRVMDN3XhCMBQG+W
wY0uDo1cHDqv2vixuDhmRy3V79Flsg9Z6xVJZ4fcyQDOllNnXKBnrzs3iew9e6K2DsnbnlU0LhrF
2pV9bBN9VLBi5Nb6Llc6pOAJlY64xmegqqX/LRXCH+ZwZU5ORvVok7uaCXX6BmoWsAfb2aPT31wc
rtpkf8PxUK1zknZ9R23WDMlwXSUc6Rp5ByYZRcIvpw9eTQcEdYckdAWyThQBE3IrZvURfzC+dsNO
9tzxAljPSKcW0AFuwmCzZuwPzFlcUXSlb4iuysZCjc4d7EHRCnKdJXXDJmny967jDSgTcOP+mQEx
g185a7avVSUnpQxGXZa5n64ZBzdTySxznwc4dh8yTwHidx8z5kAil2hNibsjizdMunk6VkuogWjq
JVsg1bG+oZSok3gyWqgKEOKKf/6fI0K9UPV+uZVsgGne3Aliql7MKXBr4PEbYXSxMOfGPnNVZsfP
RHdh2Q/H3+RmuDIVx+ENfHi16un+5SjdpqartpIn9QgCZ+GfjinaVnTo3nR1rViBL77pLzuc2XYo
NVvN/+SGLVH+M2+pYu7tR3/O6Gw9CmpmXfwqFsShxgIeYMKJWn9oMR74UmH/4n8mwxQYIpwhLL3i
OLZWXJhJfmWKS5Kjm+h4RTHhYp3TLfRSBasYYSxFdFRq+FLxeo4yUOEnyiUSF0OjqBM+YIjHw/Ur
2qgZD8PwlJBgQI/XteonQeFBRXiimlRuFTvqhcsluw4Tu7VgzfFeKNZteyL79A/tmo6KdEqMK/xW
JTGy7B/pkEbZpbrVO4pfGuW77Yx+j0nYfF1HdQW9dM54FKGPoU0PvYUJtx4ns5Vdl76e5ISP/fDe
ADJ9syd30A0q5/+vtgo5D0qGuSP84eagAkULESmUIRH/JPHI59wInNY9Xf8IcpTVEo9zHPV3clWo
KPw/nlPD/Fi3V3IvUW7NfiUF5YJIwP0ALGFN4dkZi9jFMppgt0STTFuc84Kd+1l/QbIykw39u2oz
+1j0uYiOXefz0lygN56jQ+2ub8MA3WJnaEvngdDi5et6ORrgBL2wULPoyOZSyCkWhZ9NR9Pd+xlL
EyvuxliF04pH+QH7zYqf6Si2PkEseT4T0jvsNihfJ6rBp72iu6tlUV2RRJutzcGCp9sbhFefM4Vt
YKNuDsPAYiYFgSQ5zEX0cIOPIRCfxbxDSsn3AysdTI33W8zylmftkF3VeGKdW4MT452Kl54SqORX
vtYdE8z7VPbFqKH2jjzNrQ3yfdCmTGR+h1Gt65g2nviocPKBNbymdBWnkkbZBR7hTWwNg8LSlTtP
te2BysGzYeuEylXbykoZDA+VaSywuEHq08tAYZlgdWEbtLUzYPef1U/ad1vYRO624DVc87y62yCZ
Y6ggqFbdnVpUktpjCf3/1148N7qJfq+NsYMFdGeNvFJU0YlZsGE9Z2Sm03QCvs4v09JwhwqaUExh
M2V0MKHbmSzXylSzJmB0RgEZzvPf1Qf2GK0xYJLmXbcakLFomYikQT3yo3jolN9UmT8MOu8tdgYg
kDh3lR0l4rj8DW/yW5f73mA1ZRWKHbuwoF5SnQhuzvaV7fI7c4+tcAjcAwrerXOO/fwWhwhFWWus
7QE7ZDFcBC8H45HEbKPdOsoAXDnUSpkjTBaEsQTTdFtQyVN41mrimk6Q1+h4cezoQ+LKXknMK/hK
VSFE9BFzr9ydkf9yebdhsjGmVzQWNa5D7QB2VuRJ5w47G4lTWdQP7+XmbT5UVlo2t2/YmGqHaykZ
4RbN4ktoFmgGZkvAou8lSjOTyFoi8u4VVUXB1TGLShZUbxz8KdV+h3EBampD7GQwj5p3ByOxs60Z
pHAkvGz0WC5NSha9KRysQBX8TZ1fk7ufKmo+Nsrbi9YTSu190/t032btQ4OJV6qWUIKWYXwuH6bi
JUeR6JYnmUMSUlaVghKEkdTz7S8zzl1gyQgHlIzXMM2kRwhBdT0g9K6SqvWjnf+Xxuudo0/1w8pz
Hwkp1RHJ1sYd2hi1Omc+hZ2ANdvn8Pvh65paEJmj9IuxCvxhATPGS6zlVjv7hp+wKt4o19OkA/wp
eq9ZPCtKgmqhnXuVrg6Zt3opn4p7ur03V4mXNerDukkXRhOS6/dZztEmJCoEUNW9K3lYhSh4Vj7X
gWPg2j+bOeP5D3tZ1uGOONT/OHGhijTH9zYFoKdQC3pLmxupWLx8hG8TxxErcQmB0v6mObMXLK9v
YNLJmDz8G2EItBllnd1+NBwn8j9Uiv1oI71OtEtYyqp6XB3EhO+h/VDwTjhRf3fJ13ad+2dSiLzn
1gduJiVFu0NrWFIdhwQGSMdNq7u/xY4hMi+ItGVAbWMN5jPhpqShbPD0sjkIdpw4KgZqZTqzHchS
5phmQLyv6KsgfnA9pj0sqGCbkzLPNggmX1MIEOks4egk1j7ouL0fBuanLxCzRHvGshQ0+lBQFPe3
JV+/b6Mkiba1+bS2X24Q11i6z69Mn8rfAXLsoCD6rHfJwQFtrDDkj4y41DIaU/9Qff/YIlj/W+Op
vFbcVBBdb4nefz/HfxJqLKqlgdvW1h2j+66psVYffQc4IPyTVp+HwglbO90WoLfsWtB76xJAwcLe
qXv9+NsywmveN7Z1/L0AKxeuvYdIWWFuWeZCKiBzMdMUFiyQLtM5xo/tO6ba/bYINpVR1/a3vYoG
EuOoBkAq3m7ON8FPb592BSq3hnXyuuJinsxLUoJBSwo92Rc3Dtck4ErMczUSLsoHjbUM3TKd0ddV
NQ5csXXTsFzQrODkbrukRo3gJVYOyD9Q0nWvuttWtu1EdeR164/9C5j6+AUYbGZGv2pbPaGSESln
LooxTyPGNug+HUplfWEngxp7ihFyyCZUT0avVUFJZuh7XRSeC1Y9i19X7o2QrKexfkptaB+oXTUP
wpjP+S4ZpXt9dLKHamPaqkKhQhpzVckuLvK8XnzkTVpRYVNbbbMRFH1N8T1eJ2JtbM+7W65Um9T6
P5f8mWrZvhJV4/BC7r7i3jTGrlTMTiF4OsooL+ZT1qKeg/Bu7ZJkuBAl/wJjyVbEgWGQdpEraTvJ
mRsiNOKHUhatx15QGTX47yWFRMyPnFNGhvqVIX+x8AmEA15nu805gJWhvKnBU62UTO7QCwAE/VAU
nQ7MILWTzg1ix9NBMl565mTlL1r5lDlIXbnXcnesqCwmsijRIJ10ONLrrStYopA7RsTJHfQNRTsk
jZaqNBo/5Xv5WqPhlFrQyI6fRfGveIxjwtnQX+Vr3oT6Z8fVBAe6LREzNakgMjFnxjLF6oU9JZea
SyQJpn3fmkR3PBTVZwjQqgwNypEIILVGejgW6Am1rvJWTe9n/qIhQDqiLnzI+HF1dh0gWk3YNgIe
k13KNFSp+U28w0rEol4RNUBrERWphb13SpffNNHe/hto20W/NHIXXXcUa/wcaIefI4Nto4m6inoF
CbmFU/6mb6eQ6P5YpB/+0aUVzmJ9jwslHLPHS2DgkfwoblDeVPkSJ23AjPaw1/zTWVpLSrj74PDW
sj0RLAVHx/6CZP9I4ggwBf1k+IkPihotUEyrJtlh/N2kbn5k4qlBCTuurynMEtu0Po/WplX48MPV
C2XilQjWZkBfGfdxSNN3GMJdabkCfJ5JuFvdCotYMoAISLV3N4kDxfngl+OxJReolBaeWEuHijpm
EeMQXybZwVjDufm66OIxzS5hsNhVaNR+SS1fKuudCi51DpHOKmiWVtbzuSyAzs2t/KC9wnBueVdB
ER0OFuUKfoT7Z3HHJppSh3+c9Mv6lrcLzlyeJdyXtEWvWMf+gsWmFiiq65NAl0tSuy482DLBWifx
HOYTImRUb5NLA8OeYonIUiqbK10/hSuV4mX4hqisp6ZNo09Uq4n4glaCDcHqnqGQ42SRq0Fho6Gh
2cjrAi2qzYf0Yy1SSQTOToweJXJrcv/91KCRfDAK4J6RrfN2nti73Qlfzc9gb2D2I7/3YTFNTFdj
VfZ6SsAJlWi5HreMGE3RxCjOkly8yiMLM+Vhpfn13a76fJGqaPLIC8lKlaABoibib79e/0t5SQoa
gZMN3To0dRJn2JpF2sTCw54TqmNCsNyuxlNZS5fxOK7XWyuSuxjlip0f98i6xVhoawykZu4sGDww
/8d3NL/oBzLQpqzL3k/j8theSSnPvzjfFbJwd9S3En75ZnJzK9Otb00JydGNdZBWrYqKNQpwob/p
kM+zOo5E+AMwie1KO9qZ76iEe0zmeHqIMn6266+BAvDyYr9FmRYspcKtRCd8ewzQ8x4LOrCR4phK
Lfauf/I91VIgkJ4mDwsANiw7bN+tkPxnCGSAiTCbe6bUhGRmqSVZfJ7ZR0myoj+cMeHANxcWjaws
tWAVOLCDRSNVj/XZs84mVltxU0xibV1S29wcfgpuCiUE85DXhDhp2Lvt03Dm7GG7VtI4NsF3EDIA
Wf78GAfv4fMxU/275o5GBM/pGa45MY19NGGypjvw1h9TIHBegCF135AW+IrVqxRV3S6fL1PydeHQ
YokvZWFUoXEhtLFStxrcKIdq9OF2Zwa2Nt+W/ISSfDemUU+qGB88UL/o01BShUmu492y01zIFBl1
pz6X+GBvUR/Pqp+7gYVhQsSWlx66muBk3ZCJhoGjJsY54RI1BokQOI38RiehzETgeCy/eVrU2sPZ
S8VwmizS+kgpVuPqzBGfXKSC9mwdLU3PNnQ1Nyo9dTY1FZ/JGrwa6twhN5E+9smdWtILn0huNf/Q
V/QooL6C5ga3a3o9va25CRxw+2QLVtQh2qdQtZwRv/qgjWLqvzqzzhPtO50eXY+frlh912wRd/H5
FEsUgAa0vXfYXWNKZdRvD/UAwL3G4RvAYIftBf8qx0Fm+hzpqhzC0NIEhC0Xltcyw+FFofs9mWKi
jyDTF5e+CxGV41nfvgM8/uRVYsOxpURTU08hE6if64bd9+nrLcmAb+r06q5ax0kL5ISoqgRs15iA
KVnuwxAOlLgZ7LfyhTpJluf62Dcw2x8UxzQ5Et4wWtwZMxE4ZP9+GWlWtTqUVu4L7H5Vqww0kjtA
9hIAmVREDef5r852xUCPvSrqOldyigSpY1cTo6hfKL7DtTscEJ4eYieID/+ecKmmxDyU9aS+bifM
57tvEOOhXtDDvwCtb8P3Fc2Du6o4jVAxWsztANyEoS+NAEo/L7oyeNcc2yDqm1vSO9FqqKdI8/8z
t9OnKZ6Be31dJRJmoKU3tt2Rb27IPAq05oKv3vRHb6RzSrRsoVV0kesDO1X/4ic3phdXC3prhSWB
GrsJZNKCGHhsh/1YOUlo8g/c2JTbTtbAkB9K/5xI9AI/WYe9mlN/BNh9FNOlFe8ZJb0LZMCm8m2t
bgcl9Zp/5hHXeqQN6DrOxl55jN88Hz3rBLdgsBpS3P7iZTCNJIZrf+FTvObciuWzPaFAeMTD68HY
/DpMAIErIBgoMpqGnD2Y3f9mmwF6FtKyY8+TUDUfx3vXA3z2TF+a6MopS0rQMQNh+NeTCQUyCo0x
VSJ4drBbpqW7U63VOUuAuAiwgNdxwZ29KpmZZ4Ey8c+NkM9/CRurrbgD9dGLG5XuSoXjhKACk4h9
Ja2O1yUJim3udDlPVE7RkCMy8NvGWIggbI7XYkQ+DYJo7a5irV2Y4jAytUci7D0U9mGuFNHO84uU
4aioVlhtDr0krvEway80kSe+yjYlMwSJzElNsnu2vF+LEEZ13RdEdR8wFJX/SBJIckgGhf9Mm5wM
tFp+mu8O2JqQ5TfPcH6Rax8J9K1xPV1lrJekauchgEOx1DqTphy5BoHiOcop2/6eU+oTWHkI7c+Z
3IHcZjWxGWXw4PhvHzGn6TOkM0cReUiA/JhicBpaNH9Xpx3jHuwN7xK5h8jqe7pSq2rQGsEFk4nM
pxhOFOrRAN7MqTkmAQY19louL3cJBrkArvZrQR1e6WBtdo6mT8uv1HEj/YmVSK4DtfBdpcskgt8L
jdr6/oW2LWqOlvKv/G/b/nn8XZs6gtM0RUFJwa+Q+CFuNJL1PYsGaS7Q0nQwgHf5i0CifLQjjmPC
QZDqAPUlus0jzqvFmG6ZRp2OkbWEOdHAy/amx2/HtZIglg6zYsDE0/RHMXxQt05mXrhpnMnXTVCe
9ExSDog6GUGWdGey14YhQMew1/qi4dRb0E2l/60YCcX2fuILrOgTQ1IeXTQ5N8MeFH8Fe2tMEVuT
9TxI3ZeMKFx0TSD0AlenSlWrCzw/7nk1ZOCc1YYd4CL8v7RsKsOVFtcVz/0lMTXsJF8Fo8Evii6g
EPNJJKLStidP5RVGqXHidhJIVI6O7b2tNX/TrWw0o0FQXqSzavh6QAR97nZFsevVMBmjF2zOHvfu
BisTalZJv+oUqdcpfTfELPwPDcHZYgqVut39KhlP0L3x0sUulSJqwhPJWX3DDVS0BmFo+rc4lCOS
n0CBGL/fW+dFq+mcQedEXaL9LEbZg0w0m+8483+JcpwK/bblqgT1jxiXz8K/gu9tmpjLPtgF6YOl
Umrx3NYeWZb5Rau/VnOMb5p2bBG+WEc5aaD2ij85V7sFstdXllmmr5jTtmKAKyH1nidld0voSxuJ
xrPL8BdhLjRQCb2vjEds+dmyOqUTyHbHMPWW6uafL5Yj5rqKkYS15I6TRhWUYdVY0bQi6qn4q/cl
JNTJwM2odh6DfgkiS9jfzwQB59Yxop5Zd9ztTlWZlp9uiunJDe2f+Gilfmk4pJfPl70LioNPdf9t
jxin2Zqjdxd25wL+ktSUQ9I4a0ZmyF59GiMGmewlJ5tRmfs6aCQEgYxpUjnvPt5LfazBq0igkCxl
GWQUO6QSEum1nPF+dc48ejli33Yuh3BXe0YqGhNku6/BMyxx3D6JuD6FzzyGg+y86ISzfvBFv15C
T3TA3+IdJ89C36rA95Q+NwE/P1zV4Ga7q7vPBZtlrl8Ywyl1v7OZzP0lQL7BeJouPZO1zqvIl5Jd
k5xcZu3nlFTSWU35reg0NMHPRmeLjce6mvn1Pko2noYY7EwmeA2uhearfx0rvRh8CvnYit2KRWZZ
xd98DL5CsKnQKhtS6ZlJHLysAAw/q64pzOjtU1CNyMLT8LaJGnm0tJZpjYEnLIiuluWWt4qDmUR2
IF8dwtYc4RV5dH6dez+maSwfQR0KpBRW6N/X60IhfPtNA/4Cecy6G5sXU/velqSW//la6XJJOzFF
jhC9tr8pLvPwbxdGC6JB06lmmZVh1PFeDlp6Rr+H9fnYii/aJtqcoTVB6SLseIKFgm8YNFjcLWgg
dazpQhqUtuxL3yR5ZCwQLe7Hp0A78I1eC2Xy3/huZ03eEsYp6Qh5BkxGoFVTSGVcH7JJQGIXKNwO
R02f19PqscPl4+UnpmYYLUNHaPo5MaQo8c5qQkBguUkIYezQ7Bw5SKQrpuKm+p/Cvt7Efxkb5vzB
7+cpymY+UQl+bwpi5bTTH0v5xUbvghcDO0Rmxl90S2936+GEjScCtcKCuFy1KkeF9ckPWvsgMcIm
392kPrHLZ7vvWBzq1KFQOIkLyS+iCKR6mWvcZkafmxKr/JUqRSX49jRhGP4RcHuYEaKXZErcU8AJ
cd4qFsgq95hW9VBomKElBLUV5qDdOFI5XUx0RzrXODpsJm1fIGRrmPYEq2OMXAvpjx1oPi0HUNql
mjIHEHlGF6fGZg4RZpYwYsfL33D+053g3v69HTpodYaxMZ5L4h89/Q2SJIuTQVD0ZY/73TNexT2P
WNiFiv3DnEIwj6v3M/xfqf60zSXQ97RkbJ+EO45NN5rES6dHpKwpYQIqsgtSNXUgEpFd0OiA8qsy
PfgLReo7GYdo25d33IQF9cmabZEC+psf8WtW5UUVFzMXlEHoc69jjfcmO5V9pdD9wIK8y2Vyoqku
esn+k64UIh+Xv6ZEUOpj/tWgeVW25qacszVaZko6IjjnP/L43QFwFn72kLa1JiERTGoM3dTPB5Q1
papS4DCKN2JSm8fRHhxHDTQHpBquFshxZCTetKnRqSjRM2sZ3YUbEh4WGzxTGKNJM1HNarSpsx10
sqT9bPgAUJLkgGplOlu1KtTYjxqW/nx+dxVLPCGcTvR/rlk3kvOP1nH4h0P85jMxX/RvJYlEpE5A
4w6nKu4wb5WgQRqK/QvzSBxdMgm6wgxAovY1VaBlGYc2QL9ilfnbiKDIwRq+zIPZP0va+UopoLh9
wGPiNSM+i+22EbhtjRx1HNVr0D+KPA6wTaSHoJ0QIdEg/MXgdvenVFikYNSPe0kG8kwynufVA0nV
c+PGP1m13VCDDhPnbXEunkaVXFLMWT0Q4qrn24nmRFYuzXhYF8gfYN/6Hn3c3CqOE4L/RB0o5zqn
IQSTIDwiLKF/ia3/K4GtTjul2yRZQRl8lvVymDK6H00Y1vcAh5BrWDP4RL8Yc/PVqg4kQS+uK2KL
S999tIpvksLqDz2dfeY2ZD1zUlNnxkPC+DeQXY905thUjQNAXWukIAM0HQ2lMETVtC+xBS6kvRBC
UlpEXQz2Le3qfZnIYYbhNQUDvYWIZr5RvFvMjn1pOvt/J8oUeLq8diVD8MVDYNpZoiAYJEP43yAr
fktC83PZ6GDUVDCGemCSNnMOigKuo0qwzqPEmj7n2wkCw0zvwrpxz616Z9i5NGarX7lYGClIza4G
rtJ1Wj+3shpv1AmZ/tShIR8mPNkGoiaDQHdol3OydRFlAhZEuv+IpSDMJ7xhULvKAFfOoRGLWUJM
0Z6B1UzGi7somC022l+EcztLJtdqowZYQ+9nC7gzUjBYqpoBDhiRv3AOmf4xNhtgGum6A96QDk2J
l97xXze44/CRiisJB039c8lJ+wMjjv5aZJJWCmFNuxG77R9beRASfxum7AeDLi5H0joG0gsooPnr
+yxvG+rcqFRgwn3m4vTbE5K7HEetmCGAy4LNJDQEArkmzTVivq+ZbutEEja3MvTSsorccaOLdggL
upnQp96jmHdMqo60RRkYzCVuMEhlgBJyJc5RSzMVw05mVl8QJZjt3dtzJbrTE0GMSMgkBJ6ESxOe
lKWYTR/HKBY8vQjMGOlP6htnWrdQL5jiBUsAI/R47zLMdEIqjwu3mvsuUHMm5HBooosIuicBY+Cl
XCafFLyBdOGfNA8/wX/X9ajHlupPeACR/+RtO7oAyerVdjnRUtoTR3kH1Gx8Wk2W7BB4shVP5AOk
jBp7GRtzFuDhmXfTANu1FAdIX9TauE4EXIk2YlQuv/nrws7lVV2PsmPg4/540PcgL8uZBQ+o+qAJ
97wqdUWGiF7LtH7T4MK+dQNDVOPFA6URKt430k9rbwt7crp4dP2A1Udc3licKcz3E6kPWEVznm/3
aWYSY8CFEJroth1RfqFzZRVvGa3A8s1FejI32BCecuJgpIwq9tgFevtys9NOhUi2MZESzlE2mjWk
z+aUsWC4+4mRnsTA7sfgxmWqfaZBG1/3lM/uvY1lrWPVVX3uVBaUH0oRvCGkBwlSvceNjXsxd44h
4oncFIpKMpd2RK9MSOYKuvF1JUT3nJTAytwkUrxMBrJ+5XD5/pBFxcqBCleR109qZ0faSmBf5ULn
x59vnXRgR79Hm4gMbard1XA+JoLsz3WKdfAVrNSwAorTElnZX0O/QBm7eYRL/s9+VBUTQQ2+8otg
hMsByORh5Ia+cE4DScoXceNa3jxVqH5AjK+5bK6RUZTdRCr+oFMSOJmQENVCpWOfkcj8lPR/OiAP
TUiT/pJedoJLePgOjNVsNF1lKd3ZKgkeEmXEQRwmmRiNZFatTcS5JYUJj3+zmSUBww3M86oweTbT
e/Y9Kq/47ZR39hFkGvjNrR62LEDpa0dkDgKYeYEHp8E4IDKHne7cvAvuut12wOx3XG8vqJW8wVtA
IquRTPCAS52KBYBfGPqfp7BccVGJzIfjnyGlEV/jUkC4P6oBnic+92EjO8g4Sr8qgUO3PgBUSMtU
RbLnRzFrJ8ctu//CD7KUhfXRaOnVJZKmySCGhYxrFHBx2sqk5jPE4ZYg2RWYvvRjlFi2E7h/pYKK
+ZmXsBAfAbC+dczE995SdWbCDGavTp4WnCfhduFBMEHR6usO26UhCDF6uR7JwhHaBLLjRiqUb1sT
pt7BGNRvVkjs2eDH+bMLclXJhzYbd95DVmIfIv6yMluKxb0Vn+XpeYvMb0JyiZI79AXs+81QXhKv
12Lma4LQYdLL2KPZIEcZAnbzEWEW0t+cb13Fb6ZYPg5RnWas15LQCMpUbH+/bIUXmTmD2Rh146yb
npHK0oLDUET8wpWonfxBqLKziIdtl9LCA9dSujSDgpKqheDuYgPgaUECZzskrrGE855S21D8HsDT
+rR9AO08s+O00NrJ2q81nr7yWa+44bwAP84ZjoNfhF6BsDYb8CSSkUYwUlGGzrc3SipPxga5tpmC
WJxENMRTo2/AbcS0rcjR3VrEqJJjal+EKlhehYT26E4VZUXuu4WynWIBZQeMzmQ2lofWTpgti5yO
pDUavxUk+GjMVpEa7rwlfgRICXDX42+ba6pLw4gtORj6+lthcAKqPkbJ5lfWJNiVMH3HqCEsJnpJ
MSs4/tmLbJ2LZoVyjjlvl6kgGAXw6V2Ux5x1lDvLJjbKjPIF50/vdhcO25Z96CHRmLtK7AzYPm0P
3QV80t+ypxrzkOddnsIR480PZuF/gCS9LrTXNH2EN2KG1+OoLNHPIj7nvhL3n1X21GGa4yudpKNm
BxMULVFXof9PBJwAr3e91yuVV6rJbtQRJ3xmbwNEQQDvqAK66B3tVfpiZerYbI0f79DjQZZedOXb
mYAGsYSXIdZnv2Ss8YVSO8luqWX0lx8R9QqAeFOsnD0iKcZCiwehBJyKsRaJSwESHFQh
`pragma protect end_protected
