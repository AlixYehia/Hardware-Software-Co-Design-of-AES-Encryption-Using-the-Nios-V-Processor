`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CEhloxapnNTGJVi0O5UWn6qChs3CsUpWforGE9M7WRAG1VgD4dVLY/vOqxOJFn5w
SjNy2+vPD8dKypL1bGYnRg1g/WhZTaRlhAa1Oed9m4b49BKPmwBcx01ilR8sIcro
p7WtRlUbz/up1gpilUrznlj9MZtAr9qeuiabTwsGqEU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6976)
Bwl6KUZ9B/p4z28UOj0KZBQpFwVGqAIX7Up4YUBNkw03ARtKn6b2EF2lzjiX9lsx
YOP0qAQoByIQsqeCcF/gvNsb7HrZYmTO2ZIkezTKkRUNl5sWmZetf3ws4dfd9ShV
4cDoplCq81MCZ1tmlCGh0TEX+spdziM9s4NNulk7T50nCaqe5n7nA6yUdCVhk1sW
bva5wfDR691bBrnE9wkPUPohpAeVoP40SjmIFsl0DT2O4BCUnK8NX31dGm7+b/NE
cvMagH6D33mS1TvkHhAEoZwiCcuuVhUV8otTFTPBwfUchhWPdsimw4K3bKg3tI2K
GeoaLRjhxxjDY7i+APZa9gyYwJtO9fjSfkU4VFn9U4TV2Umcsb2nqkUKEqRdA9Rs
1UlxlrJStaeOkJdEM3kUbP21dECvqtTFLKhyAaQXcjNVl0Wyu88aTUdZbQ59X3rh
PlcoNrHaalJovfOigK94SObcn5MLHDvZHrvc0388PeKxX8qRU+FX1HS9/ABQiwU5
+b37lHGd8M4uab7AUUAeMYz3w616ZN2I3713quHOId1c2rMyhZ3TtVIdrtafOtzq
h6n3iSLFh9NOvutPV6gF/R4x7bsTJrFdfe8ZfiZnF+qHztTe/q9JH1dtfqtCP4bw
nHlsNK4/AaiB2Il5S3TrValACXrVAqpvMInq12/BT2oTtCt5YzgHK0LA98DBYGR7
WeJVs/fOD41foZQcT+v+Y5u6Mhc88HoLRsgDQvsYsmSx7KwNs06JNVt3TMOh5++G
9wEi69D5VEh/n/VQgy0esN/kkqpV9GmiIMKSQ2DQpFzgmf9yYhUw3OCUzNBCRVgX
EhkcLH+KUu5euLBjcGWues58Nj0bbaWFO6SUuR4JbU0Mz0e72Imu84CQgZRGoN9W
QHQx0mw/VG40BsABc8ooPRXU4NWbAfegr/iosduHeCavKj9wr0BGTW/a7h/XdRpn
9XGjRxAVu2vREJm8T0tggiHBNDp7pD72yqIy3c5+Rry4ZiaX6DMnCvQj9FC9VOuF
MEBHXUiRdPNLYUEQ+yqmgamVqanDHryf4zxqgvb/1LtE/Z/3819p94SqJPHCXn1n
jG6WSzpnSBaMpfr4gS35YtOmr/2shHvHJLGmfQ3OjeUF0947EA0rCLZt4SYNtuPB
ID5nNIxGKOlYr8pfcvriAMqNRbK24YSgpD8N2GXGpq76rgCGOkQHFgViinGQv2i2
sffnETGxIwMOsHYLSQzR9/kgOGb929/5cHgvwTiaSdApNhQFY3artriWsV2rAkJt
0R4iNV/HiX9hMCie5OjA0lgw55w57E3CFW5vYt4NaNgB0Z+6ZH8PTMYufIZuhL8o
/RPvEpkZ0ncchIRo2CsZfH1b/Ke2IF1ec0KZAqh2+4VJR9UUM1i38VtZxHlwV105
29RE9b5LVEYq99ZZMGJpwyC/Vcum1cvDMk3KQyxB8yQkoP+tNxbDtQfnqeqVB3N+
jsDiK0ww5DdklwGu1zKSHz/e4SXK6TwSEkwLw7BO35ySF31xdBCG2W0+BLAvPmx5
/PCW07hkkiu2iaVactcCaVJ5CgnHeEasYQFZusAj9F739rB7J0RacM7c+SaW+g4k
pzNg1C2MaYrlKalqlPWu6ZK9vLao5B6SLPSVtXDEHHnRMhUYdY7GCazywvKRqh4q
pQS6lLsKbi34m+QbRYJv8+UKlfxYq7P7OY+2xTyHjbsdTEW6u3fIgkkxHSaoBFii
v9H9jRYXEl14YGA+8Rfy6QRcAR+T0te/BVVJxZs7aPZsXgGVs9/H1Jc4k4q7swp+
lqsOdSV2Ryo+aQBRydW3O249eq/hAvOlRoc8K5MQfRWo3wsn/53M6Py+4/EP9e21
Qej3gwmdx8CGNYnLT0f463G9sNO9uvyQ6qv2Qa+Kw6e6gfgmhhCN6EmpcEvLc010
G+A8R4K90W8ELdZvjcszdCB6mOVg1XODYy/XoNyWQcHE7nBoaQYmQjCwwYCPooLB
PEm4qGYAz9jtUa8NjSsTmTsR8oIekRFwcOuKh0gZcdAO7ellzHcdGsuKL7c6YiNo
47m/XTT3fnqGgKgFReLKxL5kxSVoFRwc2IwDY0oFhLdzbls1MV8pGh4vNzRDbb9b
haR7ovlh3t3lGr8smDj+QTmTlaMnsrNee8d8I5HpvE4KOUVPhdkLUso1sxyC7EDA
gSX8hSJ1aoN/bOVQPByuyz4zZE3Q2GXRVSh1spaEkf3TeNK+fEGXYJEnxUHzGoUS
py9Pj0yUDpGeHvlwm9IlRBdtEaHXjaJ4ytcEiTSbbjATrjnIBN5LlxqALnDWtfFr
y047KAwvHuZpksy0eimQ6COPZzGIjntg+wZlSYsOq6OpPwvihZxiSHYzaOilQJvK
d7n9jzZ3WQ9QXZns1lqH22MNuCex/dOI0go2nKwRC/3CuItCGNftfeVpMXiPyWoD
ysjPUj5mkRvHHABLJjWMq9MjsxMXNxF01yBwarNSkOZEwrYqizosfHUvDUVNGe9v
TFAy8dxg0HyJ/0Dqlcxuf7wVIG93FoxmLco028lNwSHreCDhG4bSN7Aq5wXTjaKf
lv/E8D6WvLDjgpjgpy5w24Uuq1OI5e1H88vZy94cfuMdON0tKEvneroF3PQZWSl4
N9bb5QsRuwlf1bHQ9YWO/uWsATlrIpXc23ofKXHvTRdjmO1Uic5Ee9moh5CGivo6
wUIzpjeUD0Dm+YBx1PGIm/k/FAtIh4q8n1I3B3Op+9eW0rblyAjQl4orBh112EPe
1XirEqsV3RJLwnFIKyE2IzBUVz7T0K0StiRJ1RKHwevJgV12htYbiU4HUTOWT7jv
2Q8Add5Wq7i7EkfBZTZUCjdt5pCRFWkdTqZdVdXC8Mo/fJsK83a0VzPWgqjYwAJF
vD+X4ZouwXzRm17v6tIjb+MMVo/20ppYIblGZbLvj6zMC1/OUuflsD9XLm6pS3hy
yg1iF6TJZWCtu8ujHVHqhFSHRg+PEkzUXcj1e/ur5MoeCnVCHegEJWOag7IOdd6a
b52pbqDX0GCXpGyalhDBGMgkMvN8T1NzpyVXrdFCQ9GUy7mRWEde7G48d0loHQJc
S6FTicomuE67LmR2kBxj7zGk3E8ywjDAN4GOJ4hoY3iAxNPoakn33CXXYj71q+0s
Fmcmh2MgsK2aozsaYnlShSb36pOHx9jNICCB9CFm1XmEWec6hp2EssjrynNyxSoN
1uiVq/oIBXWLwq/OpIH9X55NKqDj8V72cgiOtDnwwJN52G9vmV4IkvPYhWSxQuln
u+AWl3hbOPO/c1AtN3qsZdrYXWNBhWIu8BB+4zSM0lcq3A05sq4l0R5pXDNPZIzD
JooNlaZ0ypBWVW2UfeGbLwH5x1jWYnJN91tp0wN3vF0xWBoSOWTSvBS7vcTPx33H
josHOXWXnGzNxONFMrtm68WIHAlcR+O9RYYWo7PTmxfgvqBf4AzKxQ2zQqzmMt2E
KUxUKdSOBByWc6csYtZiNOiJmOqpULwCGp+NbpelaKb8CYZq//rEYMFgEEGicE3x
Suu75NT/THG3jfxOfhX9qGjf+FULNPy0v+322WVzSxD+AOyWIy3olZDLQeTXuWoM
+z+c7u2MMram7TZCXFzZOfQvKw/usHuUmj1b4ccsrpuQnkgSMWPaPWkuJ4q3jY77
y6vdh5RSECCRqn7Iu+262TE9YW0/iHz/a6HHpeUxKwGJcQFdMHVKy6B44H/kpXTY
qo3FElr3zHfRrhAIDUTPotVFDnj7v70UTVr+YFdmyrI9L2b9UfRHBzRuCx2RiTpa
/TgeE9D1HiTPt3xZ4vHEQCA+h1X5w73b6paLXrBtrP/zI+VSufz3bQSvXnftIq5S
x8ZClXHNMA1GXbZtijln3rRGJp5gFGaVIepWuB0mCnOkNEtz0O3zMtRQgfddL86u
UifEQ/ZC0HoIbWORTESiB72l+1xAnscwAr4B6C4RWUcCn04BugrEnphYZH3VVIMA
xrWHg7PtS2pwOyPhwc6eXT51E0cvq85+dB9T58sFQ1A2K/W/5bNZ3Icymqs+Po35
RdIyxu95zo4Cpip10GkSmSMCLRkZf7O+YI/G40uNuu+7E9qygjAE2OBqfeX23kAQ
rXxsTFh+KDd8gn2D4KHboy/Jyol74erU+ERyyD0Ns3JPYs61o9OM0O3dAj6sREau
STJweoAdVj01NMrUFaMM5UbtiejBJxm+Y9jFRRs6rOQWYK/gxDisQf1eaP9JJ8p+
t9jr8oxI945STvYdBRzDbVOSE+PXZmgB5+uEkbYuk8oTwpcjjWcpFgwbie4Madeu
Nz7LOr1B8AXjlcmR/TOywCdvkpgq5CO64JvMl+LUn+g8JIs0Z/FealpdMaZXoSIH
uFwtGqgpDMe7Ncijz6LOj7E2bYN0oqvWwWy247OcTKCSePlLJyFXMWoKEnn8o88z
9hTBAtR6gP30c6sWl4P/riMrXoblegqyAwa3jQKfjenDAaYcBpUOMTc0mOllzScx
bJS+N6QxKUQ2z11Vu1930nYYvh4suAafsC2chRYV8dXOGZhCk9W7YGaKBV1dEFAN
MwuhKN3FvJJFvmt6UgjN4rREhL90GbU1KL65oz236i1IkfOpA6BdeoL2Wa003xIz
sunx2WhOIiu8sPkPHuSkxUlkHe/vOXh2qkiiRA8w1mbVp/z55ND6sdL/SPoSVDrX
7lGVur80dPnyOScXU37zj0dWilB5R84IIr5rzAOeix5vF5xR3io4O+9F2yEwzXaY
eY293hioGxs8TgABsElZnCXpUFQJx53L54k6xhLQSFBeARcTGAAUN7ZrTFrhohNI
WsSnyUD+muy8HEa8/vUAtFxY5ZAMo2iVUBY26IydbLGEV9qUohBm0a5h5AjcyHP3
dGIpTPZacs24H8ZZga6ns6T9CK3D9iqD8TKcDJksa6KM+6ZgeYi5vEr0+2ZcFsAK
8/GpgRc0ZhidpBhAscdKiM6xRQ+rNqCAd0wRaAKVVpoW27O2D+gtq9XFvDSkRKV4
ssOhDTFTAdh9NJ9qAHL00dsL2d9v5EUYHva1BQ2DoYTpMl4BJn0sl2jzeAc5lEfq
MSI4PFvjsU496RtZM77NUnSWC67/9YZd5oYhZRh4Z3iaiINIgdYPSCZY4jRWosyi
C6Pl2VQrJisY3kcbZKAn2y9xVol2n9HJr9MOzdvkwdp+xNSRxv1OI0l3ysQyGYX9
cg48MUcdMeK7+yW8VZ6rA7TiwwSbblMNL/23rQSyop3DPhuqfGUwyrox+bCargWB
jrrt9gWj7W8yA+EF0G3GOH2B/MBclcsn7/YuOr9Y5Bsbp7KJiVkC3FtsttvGZSPO
hqX2DpemncnTLEO61tZ5geTw2cmP5Yill2blMVi+P5GtDZntHvEHzuOYzplG5du2
brApPEQu5fs1xeKNgdkXqdosghcTa2wgRL4A2lNdeXgsjBFHjf4wfSKIj7ayMA/P
R87wEaA+mw1/vNmJCcMq2ennQC/G4yrFGQDmJTuldyyALo8RUhI6AO4bJ/8OZoSQ
iA3Yzg+oWUxfF68qf/lYUXdAL2tK1W0Q+7E6UjlqmeIs30O2caFZY02weungon0E
04H/JhqopCS1ut2qbomxBtrmpR24aK4puKECKwva9sQ3FAsQqvUky3MGSE86ZPkm
nsw5eD71BmuLgb8e53G5R/ELULiH/XmIzWkQlxnIrUL9PYyITcXyqKsqLuoeKs0w
A5Z1IO/THwzHBq7P9flNFFxcRJZgssrCbNC00xq5Wcd7EMhwMa/2YrXSHOOQBmo6
yp5+BII6nbZlaug2lVEHkKKGreiOuM7366fOz6mxSoFaIspf6577qdtoMQJRz8BN
jHyusKQEIwlsYvv1UlOhS4HNmKcaeyRnYWnYlyZzHSDwf+X2+DMmpUrRaRJMYNv6
2z5uegVBGygMl++NjhR7aI7SZY1+4RLQEOhQyndSwDw565zh+hI5380Kug/D6Je+
2tYlce6f7qTJbADQrFrJKkJ0BfylvJoKaVaSkf3wjUih5lW4I7xJ5NDuJdyI6dRN
KwY8dEceMmdxOm9MrgCoUsXPGJKodDCBbsVHhbl/kqDykeIaRINL/W4buQO+hVpQ
ZYhrVeUA7nrRz+pnvwyqLQ6Y4m6LaLN1IAzu+Djo0SDxIxhQ3aPiSXEwwfi73eHv
uYuLMWJGoIVXr39/YgyIEUd63ZaFLtzxHgXs8WQcxBQJWC3lSt4U+XkDIV3Hpjsz
j3qjVwCbuEYBr5trgs0A8Ki+yaBsbdHF/M0hrfVvJRr8ChxTLmjHxGmyAgvDwwP2
h0cSVNycHb8c80vqloHA+XFVYxy5yTOsxOtd3mnS3SGhAMfVPS2TeHr5zFIMVjHg
RrUy4RpskUNMtcO4TSuQ0Xel3+7GhWnBy/o23vIAkt0FYPt8ECPWP5E1V6TKvq/P
qkrLCnNA+svB6982WW/nTvotp7VtKba+Z9tYIhY2cHZze1mYqyeKxx7fZ0YpoLgE
aWwlOn6EdsFA/k5YApuSl7zcKJQPMALnLk91S83+qkJZnrzPAXzF4HgvfSQd00nU
hPAiZFo9tHjZdwNS62XmTRB51Jui75ULH+TSW0GzJGmxrgwNse0lwdoQeA8Nrfte
EjzIrfgKo4CaP0fE5KRFvw+Ab9nRQvYi89rEwiNQpCCpNmw7n4T9XZI/jPtFp1oa
PHpdNRrKr81g1ExJ7+CqzFvyLwVeShcLdtVxkryEO9SeymLqFPWjBTVtgOzZD09t
1tnWQIPumVyT0LAV1LdePw4cb8KONtKBEEiswLw1fAZRUMg6gblWrK5i2fUiQ2I8
28Ab5Qpg++Ad3sXbPngUWduybco1TfAalyvKqZY2lCXKaxnDtUTMeRJAINGyZVCi
7c4LrL1q82XgwxhF0gLcLDHq1NmDTr3A/GKLLG+U5Ov40gGzE/CwOgXWdwIzGjtF
JspAIFpLljJD2obLHE/OGST4GPw7mEU8jR4qKlUFGMsImhn22xurfrbUNNEfFzLR
h0cvNDOZXPnkj9V0ejwJff7t1DTHnsr49/Gjjvio3d0CXa2HVIx/JrXrGfyMTj2D
stJL0jFV2Rp1QfmDwmbPuVg5q2bGRna9FgkkQN0mS+sDYbm81lyiH1g3Gu54/i/A
O8rRVuSt6d8i8Fdcsh0/Bsa0A2ravKNlR4NZZodUdrsDp2YQLbGp5ld2BI6lLsWB
uXwRjdJKwlT6lcEO7oXP7iHJaTUqCsQbWmJ7iL87wvjwFV+Zgy44Xyj2jDtZpomb
6t1FwFK3ouZnmpnRA2ED0Zi4KRDzYTStfPVTcxiQdyMlxp9nf+mFDtYu/peEbGYl
fURoIyi44zjgluv3Q+GNVzVS/A9hFd/yyf1aOWL5t5G2S+iDwLFN9u8Ldmb1iXQ/
asajTh3Yu8xPpHgF7oTHyww5i8zv6hD8AeY1W2hsm5+ZFDq3jqPRbZwzdx2cPzHn
WYcH3Llh9tjAfxiYBq8f0E4M3M4azwevD5nzbRA+Resna38G0KIkF4mygnqGv90p
IUypRLHQ9iVtFhvdqc6qRlkuKdkycJoi2PJLI+eoriJ8Hw3Crm9OQU/AyTB54GQm
Dr5lVY8G4vWiMJ40E3m95qBnMO7NYQKp61+mOvc+nZO97+cBBo4Ud9r+eVe2eW6J
iEOayWpYbAtt3vwkHSG5ubrQQqvc8YyNPEuBdATcZCHeRljnco9GvHsQ17oeA4S5
w0niPLdyCujl98NmCRNRQTrbQ48d8ROo/5wSTUwIvWkphpzGWkOhwLYBsHCXZkRq
hF5Jl1Vhx/G/opMIQ9nKQ8H8l+VmDwV4+A+BLoOLjFaa+K/8PmyntrJsFpvKaIZ3
OZZyDr1+KlOX8UYs1DlSwU6viPiNUcpsLKsjKMQwTuj1N/ytBzRxjnk92IUYdUCH
U9cZ/ZRRP58vyFIU9DRvVnPbMmXbtFtpbJci0Rke6zNBj0RyUTj6bCo1Gi3K2OXE
+tSxOjrgt+V8MXZGK9vH16T9RlBN4LI4b9gsi219MnAEk1NbhtuDL1Zmohf4JTpO
ccd6i2RzKlqROyNrODyyGOsjjrBJjRE9IiOGpGeh4zsVuNobVhftief0WFByedbR
GnO7yuWWuKJsn3sBYW65g+7m9MdM8Tr6I92ngN0wC8ewvdJp9GeMyVd9HXurV/T6
QsExbpT/FHx+KCW6ZoHwHAIDO9cyNiob1r4q//h4y9G8XZFOuV/aLfLvRceX9RzW
d+ePlQ+FoGZtEcXwizyktr+X769Xtw1T+DdPPs8mOWMNQeRPLOck0EWvjBfRj0zh
gphobu1+bHTAf+lkIS+g2KM5Py07TSAuuVTmS6n++13A/G/aTyB869MVaQ1IKI5K
PdTTcHufRs32Q87y8hTNXowKawu+euWiORfemSEgfzToipzaXS1DDL3hdjsWiS1t
GGv6EPfalAdvMzNZkcsfFIrmwmpFSgMV79llz+W6/tHiQftQ/ebVi+WcVIe1hOUz
D7FA78pjUKmrnKIHjwUw8zVdlca6T1G/iC7/QukLuqilnWPGSBMIph2NDEdA+14/
t0tKrJAuUxpsgWJPEuZX2INccMInV/7WpXhIIieu3Jx/qJ4YoHOUl/DarH3J+hzB
CItlm8hvJ+JUMcCqNzfd8GyuYHpA/i8A+EtMPHzYs/9Ll4IwLq9/GoDYKCzYQeSo
1eq5kCmKu+LpgO7hVr7kSntizejI7fd0+EW6pGoPkJV/Ojf5QUFlAn4ovdqoQ7L4
Y6o4y30xL0igLbAsIWdkfr+garlf+vUawKiCGh4jTHpX74RklumhkPDy4Ylbpha9
Oar7ZHBvl1JCcmE4fn8MMaB9c4H1oE36QR301pTtMdpJa44D3oAhsOYvq2e8HmSP
fnJ0g+oW5dKWtPoRcMaTaFgZnjPGYHVqXSDIz9sL4mL0Vj2fR2vcJMnDU7zvMOdn
cf0DQpUI1kgQ8rUwLv6u8KjUV1cU3852ZQfoNumpGRr7klK80KrhSOMKLYf7I85L
6d5q5q6bW3yg7VAj4v783uGKT0kzTn3ljIyfJpN9ZjoTp7OPQJtK9rruXsHc4OrS
Ec996DA3zRwAbJGACRpr+JNwhKowjdLgIDUX735qpEmGOxJ9Vlkgf2cTggJ/1c6U
nijHG7XYPgPSwIzKoAMENipku65iruMlSHw8NBcopcgl8HqBG9xa6irqKfQPgOVD
5YYg9Kc6zwdz39lrGcfGbml23+0m77WB1/C7dG54k/ezRIQaSx4FBZVFjMmvvaiE
Ur1S7RhLCRPAxGZzRv1FOSNMq9xOjP8TbSpLSiLM0ngS93J/oKUGRSP26OUYgj8a
bJPgY2spJg4JJ5dRB7pTfQ==
`pragma protect end_protected
