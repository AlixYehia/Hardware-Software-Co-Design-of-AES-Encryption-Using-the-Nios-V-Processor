// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
aFEWaIiOucgDeUbjOl6YfIxqrBfzjstTgZ6t26jM5hqOw7PNdBDhADknBIN7d1idiqaf7oPhuz2s
d84mXljGactsP2twQE7aCUmzL8g00d8dBX2jzEJS5/F8yl7JsUSAnb225LMWNib4ZvGgq8bPj2bp
4fhUhIQgdMBxKKevOZy0zql65smdL2+cNug4n41ZuhDkGwBug5mEfGQZp0mtMXmcytIRzbZfP0sr
TGwGAMOCqga3dLzx+6e67DexqnysEfrjxf2Cdj1FjU9mixsXL5Wmpuj+PfoB5Emf8ZOE0xPGwife
OP8utemU8x+fd3nHSLwpRw6a5enqp0O4YOgaIg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3776)
uVKg853G4UUISe+QDh1wxxWFwI9bekFMgBpz3Q93yTc89hJ0u9AO9MBdhjNGYH65YrdpUMLWXacb
G0j2/fBm7TyA8Ml7wejL40QzKkaJaBGmbVkADOx0AN2UptfjxZGV6D9gxQxXMPbEd+xG0+NeqZvk
JHDQWvs9N1wEqmPu2rajXQFi0m/3Ui0idEHXwFvI4mKLf1M/Ay50lOuSCpM/GeLVjjFxUpDOhfx+
bejYfUdLTrhR/TcTBORZtTNibDRBovboYe352YvAGJiJzrWA4D2tsd6Pe5oyFtMoTkKM2CSSfuxn
lTf5d8GKlRp+Ick3BkzAoX+XlBfXNSUMFd32WyeGW88FaYZIp91wZ52eDXaYHMeIAxEcGP0SzWLP
W2h+EewnJKVr+eZqrZiOayAVTqzS7TGiDauL00BQQN3yStQ08qHo41sZHgGhLOrEfOryl/jyr+Eb
w7mnGlF9LyBZPux6o4l3y3iil3sOAGY/2Sk2wh9KJIhCcwjmMOYCX8cbCvqjM+JdlCuxJW5Vj/yu
6Hx53Q2P2PofOiosohub0hxjh3iUoCIxyJ8IuS2cY1TVTcIg27BYRt57f9lSuhkiNU9gMDmQtlko
oenyscmejFuiD1jCcO0Nv+Q2tmKaewItabQjZzx8ntPv/6nPxZNTbXbT1doJku+KH0z8ZcQUrA8g
cZ0H15jdgyX93LP4e+JSgg851d6doZh7HH3IHixjC7od1o0/eEOFEa4s6x6wASRYJWoknLI3uv8f
Tqoki+5NPmQkf7XiClcXZhG5J2vCSsthVZzprmj1CJ3mZENmooQIPq5EgfCxD7O6a6/oOObRfuvt
pKTumVCQLX2VhVBhkGBD0LMAgO4NiJIOwRe5HzBnksS/3Z6d+R2z5Wq2WdNj78YLUvxMUPLJSAHl
WeGsoT7tSwfc46tw3W/TyuOYnU5K8WBzJ/PcJrqLRxu9RobTyX6kwCFK8+mpeKUpLB9lAKmlZu8q
oSGLaZGUaiFsCeIbRKq8I83QlajFM6OnmV5i75I3kytkQX/jkhmmreldmVIBjJCP9EWykyM2ZWSz
m2zdluUcJ/VKer00dp9yTxVmIb1Lu87RQrSN2NO5cnz6hb8zNMNjcd9J65xF3iSiRAP7zjB9C+AX
vs5CVB53XzphYxM3kTdWLEXnHE+eX/kqO7rs4AUnIV2L2iPDBhLo5Bi6yUTxSVpzy0Zg10RVsuIo
qDS9IOPfXF+/RFRJ622mBydU6S49eR9KjIGAu4o2kawELPZ1ZcjdWdWpACpi5C9NgpeDnKVw9gHQ
sAIBCRVLYyewsSYWHvNSNgaXqmQISFmTVuC3Jdn39a0fv9J5h0q/i87rM33O+Mx5Z5bSZYH41AZU
LPUCLBxw6kX59pXckUhhZMxIvb6cZPYzlNCTIby8aRAaMrsZaKfyUUkO7hhgU1bNPdkcY8Zt7xbO
NCTvLK8eEFImI3lbcGjVfsPQapyomzcAkErhBw8A7xpj1wvyswuNhTFtymSBnmxvDF55is6gGgUr
JfmEA5RVxZ6FXeJqqHFaOaMpSGab4SvYedGlEtmmOQ6ACyy4gF9IfI56Jqob8c/ZIWYlrzslLhIW
Cy7mboyzDd2oE10SIuOSBRjJHxnOxaJne4o0FeQIhOrd+O3K7FK85r5GUW0/t/oz1XRpcrzPLuNg
850P5tCZ4s1IBYMayjVQ1479K2u4AGwfaoTJovhiOTf7UaAdhmLqMx8V6OlmkxHyivNAynSQWcyN
GA1SY2jay/iI8xaWG9Wv3bS/8KOGtrRKfaYddL4hMJo4ZiecyZFtt8eNNZ/ZdHO0l5ak10AShpiB
d0Pj2lbi1SkmKvkw+m3z1iJHt7Auy82aZRFeWcCB49njU0zFlKJfLaWeux1uTQsnEk4yt7XzZ426
07G6vl5ZOt3MKLh2AvdYqe7WedV22NsLl/DsyU2rM7BzDdzAya5/vq4BZDNCAgu3lqMkNek9XQ/p
KRYEgso46rgfZnqMyVDtG0xLmpa8mAr0+pgCHyZRYgh4Fe5/k7CSDxnlkKpqEfQREfpOtfpVdUSe
jzr6DmX0tSvTX0or39ugH9TQFlCgw7aMVIDOhn4VJpPy+ue4kccltTK53+Un1fsHkfcIeOOnaSYG
3qi3X4NoTQr6O7pbU47dQjdbcXFsjT1H2a33CuUwl7pL/iAoX3tKwU3Ziq2lq86YK3lDAV/kxX94
A7y0/ZmsdQ6M2n/kP573at9rpTLifVwqn3+ZikvoHIjUqmjUnDC2B6X02YFj0i8pE394ThIGxuG2
nfe0v0Ru/E/BUl+DuJ1FxGxN2PR1E65NpWxO5pW6NnX3cBvt2MurmbDYLYeEv2/Q4AsiuODjNgkb
kreLhMzK+uQ3nPcTxPLVhgdLTpD0qgSjhqBe3+wqanRHStyo8FYofkyklQuIYtyO2nDUoaJgcdbA
ZlnukuDkDJZzysoOVDuxo1envmH+1UKAfaAGHUcTl04ryMAgGclyglvfxZRymLEappi/pW8kCtOe
aD1BzrxhIc0rxmowBveYsmKBKtJcbDXeEzmuFwRmkFZM29zKA+pXvf1RleB0H3DYMM5jnIFNYnkl
QEfwJsBQ+zihg3NvH+K3QyBKrGswKEcKOeW3eD8oJteh73JB456fnfA/P0O4TBVDjL4PNOq3/llQ
eEylr9LWYsrIA3Nz3POyghR/+Su7HdmvwZe/SaP6vcCDeKSOPc2CXnFMnt99RFCPaIJDKsGFwncd
PEDrmdkBvbVK6BS8q4o833ECJeaW002q4pCnxYB9i5G4wzMNzZSvZqiDuAUEy19lSwGBKikE8IQP
47R9p6b15Yg9CSOLZI8y9falDpZ8ms1QSR0yLlowkyWvlIE4CzowYEcPUJaVNpZ1rx8DGaKTSMIw
8CBVCVypz0gfLXimMqNW73w1DMsol2NsHZjCjpGueswnKbXlov/ndNe1JS9T7j2BJFDnysjLoLyQ
lNMx0qIZkXi9zxRthEm4nNKVEAs/hwqLR3SDB3oFsyBuRwq0cprvIA06X3kBjwOIuELbm2KOo8YX
59YZGHzIibaykHJ5EicyiXjsOdZkXI2jGoCtoqf8gZubqnJl85QLvBJETePI9NPu0J8I4RC6CRb3
7j4coacKo1Ch5yJz1rN8CTIh9BrM9qYBgc47v9tcG6HT0X4KQR7du6ObNEaNqnGPr3umjvhVLTM+
uHvyybESSt3jIbhkh9kGWDXH3BAyA3beyK7hRginDrSDi3kP2rJSIG/7njg7xQkBLdwCT5pt4d4v
wrPi3+QqsSx2NKaa+OZQbyohPVBWmrHDR1v3ZUoMGGqcK9W0OLlkIcYYkav7ruA7TLxG1nnncF4j
psdYp3JnYhFM2799UyeKHTyVQIQdywpRfdRD4694N1nF8UvQVb01klIin5VRG9MPQEpVd7jpg7jm
Y+mLNxHzMnc2ntCBZf7EofyZjJzi+oR7/LKIdqpZJQ44xH4PfK0Ny+29DLdiWpqsS+ObCSz3UOoC
APqN4Hagpp0/GN6VlFwjIllxd0yBZkDSrbHd5KlCzW25FpAwroVJDE4Y0yq2A2kXv+2iJjpt5MyQ
1s7fHEgMQbMS2bxkc1SeG7IpayHR/kMyTRO7GT0yua6kF8+DxLYMmHt48ZTP1XffBGUAyiWdgb7l
5+iv9F0Fu6x/cN5Oggvuxz6HRId3U+pq40id0r8v8olxcU0xQgKMig/I6JdDWV3/UY3Sr8FqrOig
wz14A/bKk9NmTDIweGQF5AJxpqsWVIr6jhJTsouEUzKK1+L9623bQWBvmR6GwWCGOihsAmJK5m/6
oD0qMGzHceDLzo8fMyLaiLirs0RDcSeJHLNkkKGHrnfm0eu+xYVMZ9K1VZFS1yGCqdFtiJHOytE7
lfvBNB09QUB/eo6IoBO11eBGT1SwkSNIAJYxSw+f4yQj+AWNfIY10uLgdCY8LyduC8d+kSqdPEjq
oR/KMZX9GSofT02hpqGMdkN79VjsOpNhXSbN19A7Z+RDMiav6lCa1wNxnW6wYRRJEgsKHT3+HvkF
qy0ryxA5TPWQDaE4eyUaxwkOFqtlkhnSCc8qzSfj4hqZdHAeycKm4v+2k0s1KFcXLW11tKay3xVQ
NX6WzLMERgm+VMxNQ8+u6gV/r5zzQhq9wsDl+wZbbtlrJd8EbkKkSYKtJtvfHpD5CVjKwFAD58gO
6Amv88YSvcmLv28mc0F34hzhRHRsZorVHVqn418fWu1pHEVp7MPZZhlAxqV9j1AVXpCGhCgXDHfA
zE8VfE6qaGUA5d6EGic+oB7w/7YGPcJ/g6cKT0fJlHQln2BxvhUyb8s2A7DePmEOSdUEAl6oflJW
1zwiShBunIvD1/mRxeLLKJPpRYv65rVrbYTHqD10Ic4AQ7oW5XPYPMb/p9gaKjAa70w6mnI8Yxtf
hsdDmGyh6BH2odVAvG/2f6i5t90ERobZ/3vR8i7DwRgueYpcp78MFuAZQgvzxov7lTgrHEnkJy6+
mWo2jSXvhAlqc5h7SMKcy0/pP1XUq7wWoVwUPmMJZzC6MwBsQs3rdJOJZgsIye6Fb6MzwatSNYJc
EFQr8ZDcF3oQAAgnKeUotUwe4H6LnYyDc4q/t7A4Rn1bpzOjEDMhMuJyynYOcMyAItoFk21ZoJu8
/IygMZ/IC3LhDFtMkgQmLO4Qb995DHQ8dLJaFIY3nT1/fuTGwbPNioHg4XTPTpMG3WeOZfGHq0RJ
Cth3WN7YUo2GIFtLPGaY4OfD2+ualZVV+/szVnmTHymROchdoQxM2KTCRblz4dPHWCarucaUsjub
/NF1Lp+9lvHzTQtxk0hVXk69DbNIbyAoteEBzOAZVVx2a/vMl4zimbOyGhcFCPYdbN5CIcr5MCt3
LHZPPb6Gcnd6ZMeSsYdmLO5foCTnxmmyvuo6HcX8IA3dlVirV16WqwaF/kmq3P7WOHqwWPMAzbfY
fv6lfd1r0e6CnDxQ/x1w8F1DDEzRopV34v+vMSaare1GATFYeRwbwYF+Kjjp4CiTiDOrP5DwXZZe
pWV+uXMVpwZ2CmfVp3o=
`pragma protect end_protected
