// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
kc3meRehWCrgmfyPwqJiss3BMvvFPSqE4y+Te4YJzc4CbA4CXMKrvO2/46/xnF4ErDGCKaq4zu6T
P8UxLnIbjQHulrlc+i/5aaZAgZmCFmow3aziR8Cmx62KzNOdJ6QDOmXoS9l9pJ6Obf370k0gUmMU
kVwjQ05CfkK6SuVAwsTOq2JuRQrMKvippmxBcCxMZ61i2YLv4sOTg49DMYQ9UyYL/VUG6GiNZwu2
kmn1q7ZFQoFF6+RjuFj610rNFSNmaiNa623eWLFlSmPvTWFp64ejVNMliUaoRHw7o8xpOVFGflF3
CqQcSwELUZ8ioFkJ/V03K0HATQ6OAPfkLqxy1A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4256)
vmMdA4J+o9msMwWCzohV2YGhk/VKdM9FLIbKVLYwrKCttc422TnxG/MG1hGWHC/qqCFt+ERmaMQ6
+9Mh18WR5tbif1zPneinkneqB3223i13ox+0kwQn1rHcjX/ZUCu/H04pHfT57ZHOfempZz+10lbk
f+tJ+a4rCmk7uzlcn6uH0wBPAoOdLA6u4rIzYfsKJP86J2FbtabBdYaipai/o3GMW+a9KWeiMwxs
zwf+DN7+2eOEtcIahqVvs9hn9kwfQtZKwjMkIKwBQTpM7HeQx8pE826Keh8Koo6VNXBgdH4DJdR0
7Oyf2mCx+IFZUm/cAoHW3ZcQuKIh8Pugt4mwMq08eVMRjZdzBM2fFQ4TmdOuPCNPmyuUTX6+N6DY
xtSoxAVYIYgHqlkmOqWbsz0lHJNMqcTZDM2Lf//PDmJNwMu0ccF4KxNsV3cYCnOU0m9FGsjHQjH0
NkX+syjTE9rNNUGeIbs3rG8qdQYZdMusgfCflvIa7QxFfqbBJTyyYGGFYAj8DJcEOmlCglVyu+0A
cQHVXOyZYtXOLt5yuDj7b0emCYFSskCYgwZ1zxG+2L7G6TTaymzTlEJUmqFu1NEsFaGHxmh0JLcf
WzRqO7qv0mAPtA1p/znA/hdL2U90PwL3XB5sZrt1acvSfLGCwoLqiFVY7J6sC+5VNAyyiwYmn0KX
xdZukERsReQ9OqyQ6rsuydh3698HbnRAYXQZHu8bTO1k8kdQEgWpvYeBt33iVSF2GIoDyQzB5W4E
bqtLERaZwH+Zn7pUl3trp44ylG33QTdqYVDN5LL5ycksGH4JIT6yYvQTct3NsuUSoVHhUtFlRqlt
Qx6USeuSPROxAle0NdUp0wGBjc/yeUiP4jLJ+IwuOXFMQh/W+OY/JZ1Mx+BQvghSnP3/ZwSlEoK1
llWE8Q/ulbmRLmd3lFyDcgr7LXqd0DpXmh1EFrR6stVAfdOV+wU0qf/DeHTFPPwYmKJi+xmsGWnu
aICE0Q4mhFxgZxAVJknLOd5nByrz+mRNqkkQ5Ptk+eTh7fgUDYNgykC11OqmhwMxY1PXRRIDfnzN
6bbxjFKK6QUF0sZpc0Iw9Q2DX6WsOlogJ++Kxq4dlALpb/CJSlCC6sE5e8cKT6gRENG4x6KuhZAk
aPQd9mN1TCLjnV5lNk4S93s76NE3McvYK8LkkAktLEB6qokmbnsm25kNIyD1PkZt3slvY3LR9z+f
r9W10QUIMJspKinu1M+d8bPDXfR7TICQOAaEDGiVLRRKNAxeyNXqnxFvyJPQul7CX50ySQvvwQF5
eaE42D/URdr6dvTzpxeOHQfAX9s3l4x0N22N77SHAwxpgVVzpEdkl9KwqoBCMWY5st7iHbSz+3tn
ecXuFZo8Hs/u+3wxubCAGTPGHaTyTnmV6TBG3t7/gYkdVVilbxP0Do6lVXMyPxMy4DB7/LAbP9X2
zC/TfwSo1L0DiP2VaOZWS760AoZHQFK20GHjz3U/5aQmYYUxuzAsLvpWK3f88Bxu5u3Q6R4fuOzA
nXPjeqv1pCQZ2yrq12e0lhHVmWlLts1xizrq6sUJCj6wFfdsEVNzY56DUSVbb9lNnesnvt1+hfrz
2/iA+dgBIAvEhkoIKdWvhtoo3SrJUfYINBqfBSPV2vs3eRfqbP+72Ffh3qZpe5hfrjeDmiChpgPR
T9XpbT1GkQBoS1yAHpbqmFiNkVMS7s/pVl5w3tyCaOBGhUN7dCbzDzJjoplfV/ImDVnamDczSx2w
oVlS8EmUdnVoAISrjs2UZMbk0/psZFBhXpgQNJoqr1eGx29Z0xfphJ/KRHYyOBbocSSmLvENUN70
M3nGN7d3Rf6M1WlNWtry2Q1fcbQWdEXEaj/tno2CKdiHwJqa9bU9kc1L6nPx/fWKMK7v4cxljmfe
aewalCuasXpLhq7RAJgb8UwxRx9EOoiJ7YHv15r4nCwe3BS6xz2aGs1FZSeWt5j/UcFmvRxJHdKe
9cikLlkOiEaCTc3fqhNUlHctHiII/ixjXLeZXOJNcCkF+e4vtKvVtt2kPHQ1aSuSN4ATz9CtomyR
E2e/no6VaDq0f4OtgXahkp5F07rlJDe0UqQcLEM640XzN9pvcrtdpzhBwnCA5A+8zurokoDIQQNE
IywDbRoih9qnBMfbaLaJj9rjzxiYYKTRHTDf1orCXlH/KIGUJeoyL6EbJDD5nI/kdOVhPqr86XGu
62R/W7JcNLQHy6WcyQ0X24h4NpWXGeaK82QMeSGk18pbB7pshbnB4in6lcuLXqbqFxgjA5reaI1q
McJ6O/FF6YM00WN2ZEO3pHJTcN6JQpox76dchyCyQ+YZwmd2MZwIQIpyCwOZnfTyPtYltHdoA+fC
14ZNdYcdgMiwfSYa3VuhP1n7L8kp5nybRuOH0LCDhOpbXA/0dvSMvTJEvdU9KIXtecF6fC4fvDgD
pTFcXXzkEsMwsVlPMxrkyQKInfncQ3oKsuXZ57/HnD+b+rup4vpgejhR8Od5M1SMAruRvhwjHUKf
OaYfWC2H8LtJCQtEQP9nAAZ1z91dowXhA7hIUmdRBuhxr4KIiX5IkSiH62jRYy7GkNv+qf1EvrN7
B3/rDzYtqjy9yWuEbz93ldZo3r3yqnM6fqpHmfCM43SDESB7XYW2ZTz+XdNyT4Qnrk47LCSSQWzp
XB0astJjDPmatrghEILRmCr6bqableaTCGq1P8YLU3vxwy6IBU1qcltkQYd1SSJXeND2IqCh8Dwn
OSkSu+f/etW+Hph9zhxPMgb44WOSrRlJao3QqdF3xIF4y2pL7K3mJC4lNZX7ZSozWEs7HmtpREif
svsY4HsVr/9I5uX+FNYPt7KlLYL6IqDbihYkcAZmS7QvCF6j1v0dBXFFJjUw/SIfCux47NHrBZgt
WKspfpKkNzHPFta/JHi66oE/i7xUZHMAgUo+aMKeSkygDBQ5oAyiEw+0y4r4aLK5XEw70i1NSa18
CEgja3HNUrTzDcadQSug0omQuvmcWf5pX9GcVgA7OX0gWupYsl6h7F022qe3NjyurDE4ocGvDVl+
VcnORcl8WVrPXWdMPLc8WBgdZtnGKo+rLzUAndtHodzU/JbE4E85UJIAKsCKuHogDtdm3Ys1pwy5
/dwRydo+ladgLCbGiJVmA9wzb69MpEhxcL4u/QAnROgdcy3Uftbj6jYcBzeBol7lZFy80s6Dt4FQ
sq7DBaYHvjI4DIJIGzJDYOHCVkVk5f6fygCm7wGFuPbzNH/6R1LNh32+/eHo6bR4p6GBdldtM5Of
inHjZf3TVxkkhw1no/B3zwFzOX7kYzcFxsTCDJlgk0Tdq+9CEqh5N71l2rGgL6FAwG6LQBmOLCFY
IAPU7ZGhgeldmB+hyNiRjX1Fx48rwENLGVUdVGhEAff4Q6OesNNqJ+7cjYxurbxYudGZediY1xTT
jiEi7mwCjmLFeZW7sOvCo2CL1K22ChESCAoNgkvCpveUNCYdTxR6+ffkXYmZSGaQjtAhZ6brGqRu
2FSOY1DZIdfquMKvGaBoJMhY7BB7uCnE6p4zQ7Ek1Fc2lifbnC0yohUagNvw2rDHGbP9xKUWfdCj
Q75Ui8sJH8M9SV4/VOxlMbCo8k40KOT6UZac0cgY/aBNerOnrGIdwgZQfOztGxf9qOkwyhlwUCGM
Qk0cffTo7RoJZ/JyVZ4EXU1resUQQfgboStX+gRJQ64oMEUpT9NGcrZ+yjOToYJzvXpD96XmUcVm
z2Zj4SYB5m1TXj5WvsZ11n89TDJqFLDj5fTl4RaMMKwGSqvilhIfPmz3L8mcsuz0rze/uHTOC897
MrN/O50VLHqKniBLwjKURP+ex2oBEDVxxUZAjqZlBRguRQEAN/hQ+PIozG96H2XHRgEGSAd1L9ZN
o+bEaEqg7GaLXhJac2uYQpo/JupHYVFlh8Hs3/HE78+YKe1a/EVDluYxJP91c29fKY5y7+4t6KG3
zQw072viWGlpPurN0zYLOjrCQs/y1v8sbqEjLDfFW/KzrWMUeSTMn2SJzEtoZwadaApF3cwOXtzi
3sBNska35o+G4R2khtmRRVTrs1VhMNB99JDLmzHvhqHG5pAXAtMM89UTrHIWSx3vzrDczgWTZxRb
bS8kUY9HyIRU9XmooP3iJl3TcaJw1nwZolfspJ6xILh4WCgK2xsBYVfP60vmUkIxK3CoDnSZDyTR
zd/QlDT1TRaGdqOEMfgssDXdkbiWHjP5jYntnxWwdsBZjOpFg+l1SC898NSyummDQC+0RN1Cugdk
ep0gQ0t9MIG3Dxr6d4Pp61BEf3uplzy1VKISMVpoBvCtKzntnIqKQ2k22C7efSbYptY700JEfeh9
UCCMWsxWPJaePqxXr9JH5GpernWGmWmZKmN6DC7G/Mik7VE7tBOgwoB6MhdOqWl+PWUWu6SbPF3J
WzjdVeDY9ozUWRXy9aXf28iTXGEULAzmQKNPJcvvm2fl2pNjId6lnO0R5zJKVbzDSNDOV5K73lkU
q110SNqZmrC3ioFJ6iqJifwbLd9rrsJW/S09kwEyyq27opjWayLHUHTn1dcSkGKj9nSsUlf/DZnp
A1LGAcz99cUfFeNnJjFG7DHWwQ2jpyebWR4TDr/44vIcVwz/EMs8R+Yki4QCHq0ymorXlbSRJBqc
3RgTog0PmD7VP7xC+Lvag5HoDTZTk9C7Dch9qb8djJCIfYaXRC9gEDXMQfrQ7T+MuPdDKJl69UYo
Lkgu3KHtc/0JZlt5kGznDoh06z2uiRcC0WdnL9k3BRy0BGwOMnYzc7zBQyTnbQyD9kCgOsjaXn8N
+bIiA6e2T9mBOJIrde6+NB2RVIo85aEwKZCqGOBYosdDGLQY/m7K+AzQDEHKFp5mKl+ZwlbNq9IO
X57ocV0YP0BELe3UXgvCRfEFjlnRExYPgYCBRWww03RqvKX/Ul/NhdxUlPNvuxZy9G4D6zZ3LQko
KANSgAdPvjzmf5AEI+lTdGcBsz0AeseQ41a3ktClS+cbvfCPOSS1B1023hUGa0UxhsfY8b4hmohq
exxxDe/7EoztaURbw7TIpF+h92GvSqaoQei7NPh7Pw6NQd+gxv1GItSToDT8FCRSdi2lotC6MCyC
eIBnxhG0rH+u+5Eswc2wY0zGuVMghQBCjrp3gRyUmWa1KY5mGPtipZ5V26ECAzQFKOIWdZVGB5rC
jIwgtyrOlSe6gmO+36I/CL1X5mUZNfW0ntkUQMPiHbuHjB6xtHNzpJadnkMuN0/wyQ8HdtSobaI0
OG/4AVDNTTUsww3dMYgMVNI9PMA/Mc1w3nKZoqTjlzBoNTKCDCS+ytCAza+4WLnts8nbkHTKWP3F
E//tF3dojpj3FlFWmEJ0B13futDhcXr4dEl1KnUoZ+GBi5/ULBP3cFvNb31NimfYGz8qyUt6wx53
sCoEvE1FLNGlIDcB2bswraELBESxxOXT6nL3/Gi/ZKG27yX6InV74wouwQS2eb+kzB4CIqSd6Xnh
0WZ0/S2i16VRX0JMjZ7meFrs8m32g48+i2j7OQ+hwmppthqj7dc0t8rMVETmI8NEl8NUwmbQvG5q
+8xmxv39S/wGfBe/MuH0pkPOGs7q/dEf9M3huRLHfABF9Jzb+cWLbfMt9CY4IQh7h9StUcaEMFv5
+imHFcxMZth5OA4irKrGfnZy17090IYtgZMmylWSszMBZ0R92bQ=
`pragma protect end_protected
