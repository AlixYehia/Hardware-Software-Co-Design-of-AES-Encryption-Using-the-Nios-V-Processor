`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k42LqRPuM1CV6dh6vXiIZggYVMxt7OVpb+Dq287kpeLBWGsIniK+v3Lj4+BH8Ge/
d6rOnbCd/WLExybb3K36WhzKeK57RPTU/6rsyFmLh43XI70X5oUJrjdpqBuS+DCy
XuBcdzjWm5dubzzT9L/xi0PsXDyR57Mg+4adOCMUC4s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6784)
TC/CxoSmdvoTNPwZ0ECgddT2GgjC0/NSAn7LJY3qXAVus0jKuAgYxVavSdZK8QoY
A4XoDVilt5WjuUmizsy9KKmr1ycq5/9Vbl4aEQbbLPdu/O/LYsl35qL5TWBNzfis
BZS5Qd8qIjQt6NC818VzKau+3SW/lULlX0ef2XppGVhddGYfKL0aNjUX36oC4r5m
RNSCt71XrO7t7+gGWvyEJkewamW7ENIn78DugAXWNiYh6HjIJ7OnXnP3iTailnhv
90TFAuXP/QjhzUaXhwq6jBbVLge6ogadOFaUbriA6ikUrU+74tLg2rnpxMwmExP2
A077nBUW+FzeFNcOEPLLYPJEeMHAviRHbfiIWbIFiBvdSaCQNJTGnJsdFVhAdz1k
B5I2+bMxADp/coU2KpaGfSyeOLcusUeShVA5XPEHv7WVsObt6dGu2tcsjgIsPSxi
4PPacrl03QmTsY+0vsMzQ6e4DjMcyIeKKji/mvTS7kt2nSPuuML2vN+mXnj2wCTk
F72WhyOFUQcGA6SN0ZSFwtjGX7C+JfOLPamzXEHR6xF+LXRS538XBXxfbZxYfbIx
dXxlMNtx2kYUHk9YFWyCrFK/HVkiBUYhcApr2AY6bqqOgXIIMxhxJikrkjzzLM2s
U3t+ARna/oIRQCXWiHRRuPqW+BLQDah8f54eHI46mUoxtb3UTRNvZrvXjgfnFhz1
Nd8YMD0Gu7plJ47gkhvJiByVu0g10Q6DV+fAIhMFioMkGJG0dyKxBdiPoEEqDV/s
+36mMxdPbxq+LrjbaIizhF1JBt51HmBXI1qhqKw4qC+mbehtMnQQ9olKSt6y9YtS
ZXO1Rz5qhYVDT7yjBkzybWhq7IH2rSi4oDad0R1BFGCHsR/lthwYvnojc37w5t3K
YrHaBhLbBRbhZP3exBFO4bLZbLoda0LNkX3fI5SgUA+ur69VE0Mu/B9iCLWR5dVq
jMOpz4UHH3GfSXzKzVlW/9c2iFdAFyBWKUeQEnkzWz6DMNiIZTcfLLcfYbUZGI3O
65aTB2fERoHDXnPtrv86u+bOCy6RP7xD9mdxBUu/ClFS9OsoHtbx/0WsnoWUWV1i
8M3+oq6IIyhCja6WtQVEV3rvjYahUrpID6ZsFDRB0JD1A/JIWuX/hyP5ECLb+Tu6
Fow0QYkb7IaAPaLvDmxgMIhMPtA9CBhbCphJXGvG/2L6sMle2LO/JvTkH/EYpdCc
aQVFlCuzxhPpe3dy2Y5CtNm08QBjH5nxSJPyNApsGfx71gCJLZ1tC0b99anv4imG
OtKKDV78TJnhBy4GoquKXt9tzk1FXbaBMAZvgVXaDKhVkpKgHU9WH9xjCFyfD2Ty
OBSwCi/YXuvgvosW8D2FQFjRn8enBMENKmYHwAQsL4PaIJ0ZxFczbDMkqcw9fUc9
RnEAvC0HD4SgWxNADY7PBVlBAZ4qcdqYpDfrn7O1JC5TsCWS9p45zZE0Q8qqNPYd
rJXaV/FFHLOYjKS/zsuSMSKPfXc+jx4muk4pKPFJFbzVrLXvDqD9eyiiZd/Qf6BR
ZclmIDQA5Hi2vHD14LGKyHZ+Mct+wxGQEObK+vKtRyBiyhZfy8RN4rI/vRc3SqRk
Xjyaxs99go7oiuvH01xqgCznjLWuTbWitbg86uw+IkalYd35TP57Z2mDPye85OQE
01n72q+6cZgW96tr6U/TZ6hc1SDrYP/07lM0p+CTR1ebhX9W+tPmNZTiN9bPP+Qr
NnAvFjiyqwzxbNCdW7NAB3qf+rkD7c1wL/DnLNil35pzZqU3HZ0887xko9vf4MMA
yzV2td8svpbTFE2YfyMrq7XtmWh0bHrWgYWxk1H/NXTGcBXed973n+vgZDvjfxcs
Mr+ntOiTboiRPFHE5Jqx1L8AtsBhxmFruAnws2S+SN7hZzVGeLD5+dIZqLXEJMBs
Ql2HTtSLuy36LdIIrjTWd0bwxlmCZ5pOY2mBI5J3jxcVAx54trIPliIZg37r3A33
vMrpELpcXoRgPyzBzWhAWUmwJcA/fUWxgoJF5WeOP4TpwhkiTXj5lED+VTxqBBMy
ATmKiIAdkSZQYKJTkK7E4iLX6rnWfEXIQreAJxJPLm2drcLsCoGOKSjwz2KTzmxd
CSENrU7FG8wNzbw4MGx+2CeWiEStvQ1yMaPk45ScgZ5meTFE/nLmG1ESIe0/PZMx
i6iSumNuEvZJfSv5qGcvmfT2q63JM7idTDo4BPQsR0y5CyLe15fUImAJ0Rvo4laA
d0JwHHwbck8JvGczmnbzbN5o6lBoSBYUZsKMSe1qDo0TN6lSxB9DOoweviqp9I1J
0PaJSBKuBolNMhZVGrkuBK1Qy1CZ7xnhtfFZ3p9wwSQMhGKaCTVyoYhAlLzH7/0I
XBpGhXWb26vUl9yPS7cwEJzGFKKL7n+fNPOLA6xPBAONcSE2iVniu3V+eK/EaGen
UxfJyZ4X43/ylANOvnjWQZuv4tskTnpiiIqdnUjpHS6sEKwYD5sJOES3wdNEq56+
AZzC+zARfMIvF5bb2RcMViiz8cDMfuMVVUalw6j5lGiZpdhgqo6+JX+ZwQH/hrLl
S7X0TNd/vrt4vGO4mXy+gy/N9Cp7EXDiD1ngT9504WorLVz6+mvBEdMikyU5xjvL
HsNi77/BNNzTrD2F4XJaLD1SBdyuO3nv9Z9AWNnvURmUHR8XFAmr2/6gaHmz6TH/
4MwaQgapySB+EDk29GNOsNeRxT0CnfSd2h+D/F/o3Kszi75j/WYKEBJHnrHuTlyF
BLnnbMNWPEo+XeF6Jk4Lmo/Ql9aJlr++iRgdsLjg+Rd/kj6WuhciUEj3qgHjRE4m
fLY0BgX/vxckLM+7tQ45cPlzLNRk0ncquM4V1f8b0HznorWdcowYryU5WQvDqi++
i57Z/e158FRSyxwN0dlDf2smfZFfB014N0Eu4kuMQ5p17CoesVPi8eNqNfCP75g2
Q2TmNm38qX9QilIGMKITivSzmIwVBGsvgYk05HyKyCeGks6A9Q7HlOr5clHJM2jv
MJzBFkIS4LiaAY7sbhVHRIafkEsCiMi7SkZhzr23yXgZsViA+4TzHnvXWwO0EwCU
b4v3xbm029+a8unJW0aYOQfKzIoMxrdZWHXfuIlAGM9XjNcbynjnPqojVHGarMQY
vj6ugAvbyhz+tvt4G7S7zvPCW9NmGgf3hHB/s3WdhnbR70iBWB/KIu58DApLWSUc
xxdBmyqfge25NN/CR4HC6UC9dHWIOXYnO1oh9x6g57geryXUaguwzVLXpgfbBQUX
qDCloFc4lPOJuo97H8Tr7nh2ONWeb/90AOAfo0LWYs3qGrdTVUFssd4ZbRLtYJ26
zdJMmWBK6MO+yUD3ztpR9e9YRD+PcqDIb13hixsC8QiopdPfxktdzjHBM1Gv5Rz5
1va86YBi29xbht7WgsGPdewYaqOHDQSeJNYmn77ceEFHqKpKDjezvSqvz2NWrySz
nsOodUwo0TWVEYcLSBFbOWO6il8Pn3hP9xON6tWNSQkgAYZXS7U9T8YDQp+TIYoX
MkAb3HxAyX9MeqCfYpRpVor2RH8Vcf1ns3lIfVZpoRX34Vy+346kBNa6vv12DYt8
R9cjjT4rwtWGUzj5jgFv9F2NgN0tl7Fu/QBf1ZhO12YBZXQuAtwl7JVg1wPwlCls
B9d7MIOdj5tmhwaK4E6anqMLmspc8v1el5+DYYcaZqBcJQetjHVILusuyUw9nRYo
ksvsHHXaBZ5uNQ/A1T8nqRPbU1gTtkWJrUyUi9rifubWWFF6AfPLdyBlhwqAWFJv
SU9T4ou0oqyA/uf5MkvXdKwnWFAX2xZRW0N9p6RXNIlHf1JRsudVgIxXCgO7e7S/
hfhQSXo9tk0Bkf5wiho/AAcdnVY2rkt503HDqdaD4YFD6WCzRAOnELFYC0RYGcnS
6u0EAVdGN/6dt2qZQpcUH1uhtdybRKB9nvhMJyQxwR321XAMvz6ef0n/emQ6D1G4
Gleo8hGqXtPrXpyq981MKc0UzIFf/AGjAyl0hs+14NPtJKmfFCFjCf3StvgF4rOe
AHvHjWQEiLCSnk6Y5wzcBprWgeKjbzb9BmL9Vlk0jIBObnm55cPgU5VzwOyYuZ9C
JE67VTTClsq/SPN2rbBHlypWQcvdVEeMtCYIv0kwY2tG8NR03ZAiirzq7d4docfe
1Yk+MI+HnPP9rLiJEdxfSXjtnrRzkNc8TdY42Wm9YpJofSKIBwbgHepXmd+a6L+0
0XOMbSMa7VCxZdGO2UvXbtP3mpJoRWupbmo75VwoneKZVS/HYtsChp1rfSK5plxR
TC1h6ZaC1sFNVWCBrt1oKBPiz2SUn0CIJywMjsh3jymS4PkVS2oIvbjXPRXh0jyk
H+kQNJ8EnXDItsOF/hpW26AbZHhQnJzzNVJhcBX6nTD1hXlEF1a4Qki6PZmtqQFC
SDMUkWl4LcuC0X9IHZsjKqmLrG6wST40Jk4+GKsfpOV6LuvnXlEN2o9TTCi0E+SB
BDH+k5sGg6QWT7yNw9d7nFKJvFPazB/E6X9v0AkSbc4QOcW//By12LBq8P8DV6eh
brxVQgTSsnoqHDPD+75S3ppWsdIi4+FXKIwubm1keVzP9Ioi7w95o+1fN9n56gAA
dgjYocRhei/3uorQ6QxEXqimOA5CwQv6eHcvUuVH2akDLzEi7pPLm1M6ZKqysakg
Zigv4wD90j+hp0btzP2np91axoIQ+uYlkPoKiIyEOlv0hCar5JjvMq/8kVzWLAEW
Wb2tZR0kg3mDYYJxSONY+Jt3jtfHNUvSBQF8VEofaNEBvrJVFmQ0gC4yjC0Jl2hn
qj5EnRJMGNutuOPiFKNEaamOE5Cl8hzjlpx1qnQI6c2nU8GbEEk4heAcwRDoRce3
mVvmljWqagLshfWbrZ86rB6ctjoi9XXHjYK7rt2gf+mAajOvGwcN/wWx9VVw9X77
DKX2nF5ntppYnQ7Xdr7OygGA45lv0K5Ki3w+zRDBnCwLANfkWNH8hXUCkCiiyv4v
BNow/GAVlcnFLDhj3mTgJyHpjHpS5F//r2LqrGmMhaExcH1vFM6aXjIzxMGvtwVg
gp4okHbMUFVv4KJ9ZiP9Gu+6Hi5DrJRpeKUfJ/XiYUMRCg/WBwXKRdKlCgn6Mhgl
GH99UQ98XIVrg2y08naFRmENL6oBbK6prNUUHnSwdWnuckH2poxxSZInu9Q0QKBz
74u7YOifyJ8o3fCSrR3HupkR81Ape0SxjaPCCn2rSJwUL5Lon5qs4TkdhrvcqRKX
gsMKPO88ubof6TM6pSlsV5qV4HX4eTtkD2dsfnPVR3/qCAPENQvXEiLiG6KY3Q66
k3XJ/pkIy48Mbd5Rjp4W3CfJHpvZIwrgHVjFxz5++bxkQA2cAuxT92dWwEfiST5A
ixliMFpUHcYht+/x3QTOKt3xiklnWPqr75L0hVbvPzFqZYcp4K4AL19azo65T/YE
uZcvZ5mnG3acA+5zCFS9ESgtX2UobJ0IjnvF9avuBAEAh2o4qpjCmsaB8byl8yJF
LvRA8Bq8eR9LGlQzunOCwjQuU2BbNzoASRBEwOBEttM5hwUvwn/DCw3ik8VYOBdF
RO/pDLaoeKRnIkL/ELCZiilgAvahFTpWo+lKe2D5ODKDnC//QEXPY1s1AQLzNaZq
wDl8UN6J+bwb+s+7/CS9ExycmoW+q/4Vzi0C/aFgA76S4Sc/AZ6hU6irCjoLadeT
QUXJSd3LUwOnNFF1dc/I/HD6VsKPzOaMX6aM1sg4KQQwbChQkoJnZf9VoW5g6w1Y
MgSWnlNKVY5e+Hec5UVX2neyuRAI9ueFAM8sXlZnv300wqtr1gOTpi8TXcyyu212
Xwxl8FDDXhlwPBFEyUj7UE1v/COS9hQVTLTByqQUAViTEkEP3YhA1UBpOXQ+U0CV
xYFOhdVrWWE62gNc5tPWz19UHf5tI+c7tJA8YoTu5ZAs4YoEjnloctI1JreHaCkP
ROZi8IZeI1sNHL/3tP/dvjxqAXntgzqtwbkQLdhNv5Gj4lgHGXzn5NM1nC/wdBBd
9sl2/dgProOKb7CY1p8Iw2J1+sWAgyP6JRlWnImMNI2WN5JGhK5VO5Y1P5372Hhq
4KUsc/zTYGRk7nQvuzMnorxV8SG4oLXd4rHjdmEGViLe84otJ8p37YxBy+Wnq8ge
Yl5lp/IL5xz1DqyIO7nkEf/sGLAcQ9auQ0BUPYA0NzuyTQr5Yf7P+DPz5nusidME
pudR9wRHlakgWHQjHZBthkJC2u6dm+0NhKeHCyp1wpDkUoNmi3xRgJHGZuqwqPFz
2bxXmJXlVw1Aw8sDoxZAKQvCr5PUyhY8cXgT5mYAqBvzyiHCDrTgtc7Y//LubJMD
mHwMSlDqIv7IU4SvdgwAKUZBCfzfa28RYCJAPauKOrSnGCOhn+MwjYpxkJyJIhAF
H4kmPgeriPcDfMhXOhA5p5TBmtTt2rdCnTKQj3kDGcQeurpcSKlCVaheHTQh8r5j
yU2YOx1gf25F8ske9CrwLxOBSxVms8Dg0FOeAkxRL0wDXeWmWATFpl89SsMSdAV1
AM6gj8kxaYR7r6UWo+vOx7w8ntpkl8Mks1MqdjYZ66mcKpYK/BG3YIU5q7GbeVh7
a0wZpkooJzCRzr//2Rfl0abQJvt1AgzsLoHWet0Al1sDSYLLdNNh4eQuwiA5efPU
kA39uZPTWfekVmVkRoY9ciZjrA+ypXw4s28pC3TPHqRXzQfCfyytOLXSihD4cpmU
t19uFeijVf8rYsu0WalGR+FKrswl2jixJQq7vSMh7AVI/21qvB3KOH+Prc2dZnz+
Csi4hZy6AK1ilkbUFKb/YUu/tcvumsQDORicIIcs1Jb50IYO/+G+BmoxQ5n6A7HR
BffPqMNKy4EyWSYHbq6DXRIAJaR1Z+rtQ7vCOJkoa8hzNdctYy3Dj/GvpM4G3oD8
mcAuY8fJXIgKDXE7u8BseswL2V/R8bvf8xs+NJl7cDy+DY4WYhYlSybYn8KRfA4L
1jw3LOfYLz/MxxFVMk6mOOnzpGw79S1Q2l4Pnf5UFWQOZu8Y1+5FRseAGbN77+UD
UukX3S8gw2v8CRxezajPolqLkDsXqnfpVjlJEN3/ggE1vshobj+hPuQABHdxeMUT
vbKjxw2gyu5f/9mWWg2wC/ghOB+tv89cA+bMi/BZQpTylb2nxGUcid6Pa9KdRk8F
jkxGo1fRQiK8P0ofpmybbj3DtgsrltC9/+DlWjvdAyaYTkykvzRpTt54XvpUlA3C
1+ffLN5Brsvz/JlF0ESVocU4o2TUk+0pEWm67Oi5+dEobX7g/0D7PNR/Uue1VJh/
PKR9toWSf9zGpsNCk/boTCnhNYNnJMKyM04c9KUSgKInfZ94JlFo84/o7ehCWZdN
XPi68sLzyplmMnpZrLx5YvZVkMPdNaH0QuoQsSEnBuRR5em5LTdn4mcPuaQjbr7d
INQEjM+5ppg6bInNDFX4M6GwR15aXUDy6Akfr/OLmvsjg7ELjdXL58JU5hnEkzuE
5h5e1V1GVnUOthKwHzgIdZFSeCojaoCJ7enSN+vgXRv0hObofO4z+iRI+HklNpnR
ww2q56OUdbgKi7NdZaqkqFt2esYC8zmjxhpqshuIyXU2Ng8k8c4OQcfj+wdDAsHq
ZneunwwKgcIaXEPS7vWDcvlQblBXdqmsN16vzl3e+MKwMkKIOjVnF6ZCJmFkWEXu
FVv2sMQ5pMuuyMjjqapio2j2/LuTlwT4w2HPalWl/Temz9vGBVOZsweJ5Rsb6bB5
emBV4woaV43ZVpQAHcXtLB1e1IOHePvmmqSveJ188rFAJYNSJqj7WHR13UPpXZ/p
TcPFVxQVdUKkX1uKQtGVT0v24j/WUigV5J7N6SUGe6c244JvQbpyVsi6Mx8tQEsz
xLq6BZ1iN78CoRbaw/RtXubsN/GVUeuUMea2YJsmrZVgsp4NNQi0VE5c2I+nCGMW
w0w5OKvJjIKNOut+jSAb0PikGUW1jhC7h8WdZWc3uyPEHG923MmZ8ehXfm4EQErU
UewvRCzkIwT+DBwGTMEmiIaLBh9qQbsS5s09Zh1GM6SWBzd+UtIfGJMT0ueGBeAs
dBdOqz+wF844ydmNSuX+u3D5qVdHQ72di4ymzW6h2wAANiPNC0bLXiq/Y1IubOtE
XeCw18uAT8AQ4u+YNzkC8oHGq/PkGblhSFvcv6B8d0ifwQ/KgxEnMuNn8JzJ3wiN
cGU98yi1hCDCSrNQ7kus4RS3FPoQrDUXvQh3nTodUvfYTMgNNfWbKESEDDjFavLc
Z14zSK2t0gGlusucYx/7XpqLX5LKC2GlqZhnv8aBlXZH56bbEzI/YGnu6rnVMld8
Ek4vGnSjfz9Un8NRU9EJHywplmWYEjtWcBAo+Vmaiq1v6hd04x6W+zYOZ0nms0fW
ByuI8mcTyD9S0TamKNtOdPFxemFqnu3yAQ0hzkutg6GqdibgTgVynLLJfimYhB1N
amDQHAK3MJrRtacYEI741QZeLbOvg5AMP8+m5fPRY3Gjrso5newlNFdqURE7vP6n
g7fjPuatyA8uDG8TvOTGxvX1pqm8mpWQd8ZYbIGbz08LybNFb7s8h7pts3hB4d0g
94Z2zR70y0n39NI25QpA8bw4h8Ss+mKrdhBO0Qq54Ti7JzIGIrrWiygZz2wGi8jC
GOfcpzpRhJ5nRD4GBf68yp4/9RYjmbnXqhg83TuNhVOAlptM2SvG206dAs9xCGxM
sjlYYRv+4sBNtQ7CLtgTiBFc8sLaeb+oV4XgdGLNw1OOf6CeLJjsK/Kcv6USUYof
d/fG8F/T04MeWp/5/1YUniiRtY8VwLqx6XR4gWYqRYr2W6tO21CiP7ioNNzbUUNF
ffMjFMtSqqqIAkgV3oniWs0Xh3zXFrmTmW+TpQpoJc+/WUU+fwM9I+uW75DjmxBj
TKrek8GWWY3lBeFI1g7N1cJQmVciPJdpiyRPEwfMHaXiLUoFjLxudJEDmvvB3qk0
xPYhpkY1tHl2xayFKi+w+h+6tb+SOQWEhjkdsw7FDu3brVhNh39JI6lpLwShMUZq
+8JLd29hd+HLyo6HrABtGg==
`pragma protect end_protected
