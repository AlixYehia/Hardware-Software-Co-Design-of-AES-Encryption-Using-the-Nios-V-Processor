`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QaFJxHV1/lG5I+ilBEemNX37IZ8dWNCe0v/pET5Xixmr/AYLEcuo//AMMHmXu1Lb
9M77N9QPUlsMXQa6G9Mb2H4Je7H8QyMZjqJjbyuzHkESlmxfz8Zd0gwUT3TaOG1Q
kEM1JpkDm4sYcoeUrTb/k6plrWfyVtCQVxcm2QRUvyQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32288)
PF9C0FJ50rd65/j5BoMw5hSW2mKyI0DmMDiNWmjpTw4n5gxdtuldnDpQNCaw6qs0
KSq11/6AZ9KaGYzkH+RPgRCYI6C+o/0tGn1PHWmIVxf/Nw9A1a1FTJ8PWd282ihJ
SUNbOqU4/UhTA/MZymmqIDeYyFlLscPFM+tc8LMrzncRzPTyE21iBLIosYGEeFdm
Tszdtu9XNVxcm/SqCNzhFWlKcj2AZw7vlgVvp+TzQb+BjyGhhIj5EHkT7Jp2hL1s
L6sxqMGdpUeQZQoypG+1NCmZJbQQEsebtp3mNStLbsyJVmxZLcXjqqEE3OK286/b
o1BMnPYv+KcIO/fndwPGu/PD9yU2gNLzGOCx12RCP2wKY4/NkHRHd+U0F8p+QXL0
3p9t/uCnoC+wpFaBY5YfszfvPAvYrix94cVMwjfi6RaoIWKOsruE19NxaH/n7dyB
5QbOF2c7r5MBs3DZeY6D7A58E9/aTNxTRKQbbA36tdv6HUkIzfeMMqmxDCmh0yA5
S8F73To96ZTfL9hYUKFnV+x6K01T07qkvmeVkIM7kl1EjupzUpi/WJtXxKrLQQ7q
0ugZwlpV4x4MtAzW74+StkC/tfjYRDA67Ik0u8fqoPh+oLacCtYdv3iRgD3wJJkZ
BoadAw5yq/qzqL5qVMsM0nyceC1pipRAApnJAuXESZK+gfnCLrufTCrNKTBy31LX
3sL4Dj2CcdHQsssr3jNV6d6G+Be+1LN6qtj1hcQB9r0SHkuQrHn89DBvgPrnTaj+
QW9FdND5CUPzM+kXBd9tNJOGG9tiV++eZDZMGwglRDJJ5xgetX0kRbNZzOenq5Gi
V3JTBtDZHLgC/piuigw3Br9WkPYCl4DxX+OrkkPTqAJCUbhjRWRBmzRA2ei1BF8j
WdRKE8f3zjLh5YZh9AI8MQ7WeI4Emv34qCa3KUUzCmwIR6TC+cdBXeq/Il11VF5G
Tpunwfam/EAs8h5Bf6szayLKvAFetd2xka61T1qDOuOOePcdX0j7FHmnzOSyyTgE
Yu7a9dp2V7zrR4ttAFAKN5cv76CYydLGt+wedFS8ohnefGlfW41cYYqbXvldIiTY
mwrI5/HISu57AqOrc2QhDmTSXUSViqZw3ux7LYJjZf0P1LnS4wkk1yo/T6v5wwOl
tBeOAqivX19O2AYwnr8RWvE2Cui2Gh+8cxoLDE8GANgaEAVRVgHJhkDmpB57gUz6
gwpyVfCRtlKC6v3Y4fg1CbSU5jPPt0t1nnTgGc4JEFOVFy14E4YtcYhKnqklP3RK
1FUjHnD1to1puwL3A+AKBgTK84AkSSJA3VyxKoPDb31FgI/1fsonDk+9OK1OErPs
wpM4g/xJ8qddpDKvB81BHOFDORjfuPjEeJN+973BYwSyJfOo5bnVS9dvu7KZZ+SV
qvuwiTLHb0SYdg48St0LsSGncOwrmCMxYfXIkHZiKP9PByFdwuDvbiM4WHwjBJTr
E4Q7ZMwaeOJxHvcjCV63teEhNbbfpNkB3pyjiWrHhtLERxABEwCLaEtDRUiK5v6x
qdPTcvss2Ia7Ubw8XinDNhQbgGBXU2/Mr4yrIoUMQGfyRYSigO1CnDqHD8AJrDzb
yFQPnHwLbbEi1/N8x+aVXG24yzFS62CabXVF/Vc+xWYv64ugjFhE9CpwfR8Yn8It
VjZRaOBiOgouFNBb+kwZDSOeZKijssavsD0bw4LU3yscfdimgD5PXKnQ5hWV9zFI
cmIrIBDrWRK9TLMbLFtNbXsdtXP0vjiq7f7rZoaXHRqtdYuTPP5Syo9xBStIXfTS
b1oWC85bwt71kGbMeVj1JNb14R7Mo1yeJLgmY8aWny3Rdt2A6vFsRLkO8pIlxNDV
hlSwIFqxXfpcCIa3ru5d7ZTJ3b3MntlgCRnMgGfKkyLP/B7hQqBth8RL+GoFslX/
3a6iiqVdOoKrhbUsPhtJnWkHEMxBybk/RyynGY4VEQwdEbiNG4Mtngexeg9vFuJ9
7k68r8gooO9jF29Qumz0SsWaOGIgVTIc9pvWEu5OErP4LC8KiFEVQuODFQiw4UHT
biLPyCjSVmE7VrpKHQ+CyoIexUOZxEbwMLUBqkcV59bSDdxxK0VKooIXCg2+2BFP
xIFnBZFNgnCA0FjqawqJ5iSgq1GbYTGW/k9xgDYx6is9qRsvL7d9943WY2hI/WN4
5xNf/oj8DvYMU5fVhfs2NzbCeVgMd5h61WA3yAZ+LqxzudEUPgm5NXYQxacifq9W
1RxYzxrQL5HHVllQtiyRnvRKp7KazK8A0Lq4WxkrlS+xV6eJZU8YdTtsRtr43S+e
wcI33qcJki/nVwRdDv3hRbAXC1+OYFIym0fvrJ8VJXDTlwftkLsibbAcZjqxB0fn
eUaRjR3/X32+7UOl41fetfDuw0HltWFgteWDyDTz7P2v++1PdD0lZt9+akGgU5id
mm6y8O7HjaGMw8//C0J31Q2divqjFLe6gKe+NvoTCw2Y/lrH2VXsW3gMEem32WCO
0+4TpR1xRty4uJhInabUfe4CX6RlJzcxxv17BBJdNSQxamkC5rCXDiqqRbZPsip0
VQJHzS94FVxhA6w27t9TTytdIfldl7OJYuAAGlx9dRb3JacNrGbxJgKLWfreI08M
eRdN/bKR2Bg8XZkMaBy5StyFPk38ONCY6Q4THZA+1idySJONWw9MFqMbdiR6j/U6
LoABNsqFJGIcfFeCOhrbLok1eg34yEnOoLCIBg2f7S5tE8zlY8aiDHjt4B0zmAJx
1BH1DciYfwDuToA8qIMlAl2zs0l9XcvTyPd/mu8do6cLpYXBkM0HTOpHNbzm3nAF
Cv2pv3SAZu56HGIUP19Jg7+4B/Ucs51bQsQmd4Izkl0+XQy/+bth8vWdCslLbnY1
jlGnRL/hGaqfXlJTNoYpIBX869hHsjUQ0rXh0yzoSV5X67tpdDEEONf36XSwVVGJ
MLcLiSIN34LzePC3G2OYV67Ik7W3oRdnhBZpvkG1ftZd7NDdEqRvz+Oqt0pjNBzd
QzkReEoZ9M3xU90i9MSx5w7AhEph0Mos6dPXKhkoyWAOmqn6AyjvdO/zyUsQwCFY
zJYCVPZCUk64I2ZNC3IeWw0s2PfSh/XYhYiUECbPJmSTEWuxUcPN0KAFyRtN9pC7
MHAX5ouz08rLFb6jmSbQspULzPwUt2/VlLiIztGPJMR/ow3Un858kEZ/WlA1Pd57
Yx2jTjJa4vgXiZ8Yatpj6yUBdcX3CZLqSX1CZJ4oV5az0so8dzXKgOiJ9FvvszKw
LYEDizDMxd1PtAKSlKafx8gc6S6BClAWUJ16+Gtq7UmGVgagWslBDiPvbDAGW6QF
eAvrBl41PZzxukKcXxlXAHkn4JR/zxHtW1r/LXWOCmlzMbnMRV9ClQq6FnU1A4+D
LQLyooU/GtXu185RdVyjOjyyyThUWsqR4F7DywwpaHA4tFR7eyFXVrQFbH2IKygq
eju0Kgsnio4d7dcVXpGujFdGP+cij76QroFWF+Pyb6Ekqr6/UVeovicXYrY3v+qq
lNUWLdFJ1Yo9t6dNrhqIIhZd+/A8j2kPtp9XMI85m59hFoCv82S9RCO/D3K/vrwG
8d9brmvXOXtybV/IuIlRfEvzkTxUKB2RMxd5veL1Pe+FwHTP5PXOpyFS/UuL7QL7
n3/6KKOZOJuRCca2RyHNXGlhXRUF7N2ReZmUmGW+/LjR9+4mcglpHWwsCsX0HqBA
prPvbrxB/lCCgnRur2yo51QJnRBWLkWsxYP1hYEkUIEjJ+IPaigHphrqfCyYDonJ
IfipmMmXR7YKJLIQNLWYrmlC0d7iHPlUYg+vqit2rB1XGXepyN0TyPslXlUNAZE+
HSC6ndTSsKoTy51jmMDGqe5nZl3g4pRCbqam5Fa7EmIi239T9avy21dazb9FMSfw
A8b2c2GJnsZzLIhfafSU2635PtmieU0mb3Io1N1TO2FVeuedfidk8Q2CAC58CPnD
BO2eLEc/6K2Pw2ANUiyS3ZUDVkZR8RxiXPja6ZsqwScnl+/N+NKHCe751pSU5bjl
h/bDEYcjXT0LctC2cH8sPx8y2S4OdmiLbpWbnm/8U3nHt0e6oQhHfHmiCYJfVIVV
m4fST6rssfRcUwLo4TVx0pP0JLrFaJKKI6JEi2mVJcYwYfSC9mwlOE90dRapp+zK
grmBmh+3DlJmqh3WeBnJ6+kMuQQbRul86iTt7UzyyuwXfFc59OHk65LGFtgwdxTJ
OoN1nmNMpnWi1BJrelB715+QP4huz8Ou6LOcCqMyD4TSd/aPR8CBpGxeBZUk+ON0
CJNgXTxhI6u+PwEBwMztZFQG4e6cCpeaVeWYI62NItUM59ddrF/rbH+y2WNRs2Cr
DB1E5cNDnVIDXSizNWmjaody2EaAuhed63FBL0mHqIzeVRUIlM4olxuYTq7dMvxk
UY0jGm4CGqZ8VjWSt4QtSDPBNhEeDVW3w2CYbf5TbNH1zM0cRBwiU7qHmG8etlZi
DyTn6dT+myJjMXKXnhPajM2Qq+ewg8/3lTLl217bLXdwRwCJvuRWUrFpcDE4ig6E
rvXRF09e6izxodm0Ofw1cfeDbd78K6wcWwj8Z9kyn01H/wSJoprTgNuGsQtv+Kdg
Xch+0K3GQVFejuYy3OnXbMKGSEpsQK322i/MTv1jXKisdyQht38/FhyNFgP4ci8E
DO/8XReHHpGgx2fi1oSfZdMu2QFDJtyC/fVth58kEVif8sO0vLviZnSzGBmqzZ6f
aaEHusxWMO/OMTwWnDSiTQdbYEjIAS/KnOtqdA9r9XSjRbXBIoBHOCR5mlC3rl9h
GrChaMyck4Zb8j2RvhRuPVpNt9Kaicc8QSCQ8TGQ/J76NXMWb5ayrMK4hqagC5DV
cPSWsnIlov6OQReEPqnYEt8JWEn0gMTAmJO6eqLab18yFbnStpZbKGY3dx1I6fb5
5W/gSSw+wozZd9nEYs9hlwbOnzrPrs/Lfq+w/A765WAqebghFCLrrfc0rf9wsqQZ
jHo8BP7MmRyyxOrspXxJBHJGsdDL0mZUIyvX3dUqxTpD6VvMZ4YcN30d228dKG7n
qfMbCVLoH7xpKA8CGUlcKhvbKd5NUFwaXjP30eeyaaiGy2hr7YK9ZSmApSpHGHoU
oIscroQyOlpB4wI/f59c36XR3r6JRzl/1YyEoRLfDTCEq6YDEs6rn0qvQTJ+vAg5
7/Z7RNEGAi/ODMAmQgij3Yxx8p1jTAwkUSTUPFJ5BW8jm4yWAzTt0JEqnTpXP9AE
brygHrq19+n27OaPMKppee0gnz8EXZoFh33sRo0Oj0JekL1Kz7xWEQU9DhcpCi0j
ZMYZZK5OeFtoLIN8rJY/mNhGz7CZjxGbiEi9bGzxjwxT/trRMLXPhlZNa6YgvSB6
c/HYgT+Mn1M4YSr9uFN162EZN5qCp7T1WSySUBnFFisIIGefvhh1Cph4PaTFWKRQ
YeNqPc6SsE2+6FEARsPbVeiVmTR6yVNvnLyFDErmG3a3yZVknQ0cqXKWPwzokEXK
1Rp5dzxyswdW9+4hh8AC13KA7sXQOf1yaqZ1RvSJgfQ5xjXXyoL8NtWnB9OHjKP+
K3ekhKKEhZv4C2r6/ojn1vqUp3mcIeSI9tjjY33nQc7C1O3d3bimHGc+M6C7Jr2I
g6obklDs5r3WRye/Zz3suUOPmnEULm6vlk5to7FqapYYykCZajjCCpRwd8TYhgtx
oLq/XexUGXcroYS/v9Wmi1opk2CkBmlDxQv2od+dL+ZEzZjJxbeZDn/tfY+u4qUy
rKUhZ85/TOelzK97nUDGQOa/ZCpNNKbelU+1p1pwqqKjHMxuPY9wG0mE5lkFfDFf
GMa7ggAHPCaSxsNBbkBPND06kLRIT4r7DPj6l2NSbW2GBpzUWUu0MXxr77YVRLWa
pTAW5bcrP2ak4K8grBYVSplpzEx6qNl27lvVut2unIp8yxV7DlOeJdjNXJ8YDXKm
q5d/aDvfPeb3WZH9LG6GOAUXOOruLIudZj1Smhz3XIsUf0sW2RW6nAzXo1JCJmDs
Y07vah+J/wVigEICbHt8USAjZWNyhC+kqxbCdvEYrB3P2EW6ZzhgT3SNFDQp4DdC
q2C1GWKYu8gYl5+0E+ofJJxYqWIpMC6KvXLmLaNLqXuH618O9TpQxcmvLQslwtTU
NMFHlhfOq7JF9y+/Wct0gR86nxe2hp7jNznAlFLSG2/icGmnfkQf2vPBCPTZkRrS
/lmywx6egxlM/Oq3Xh1DXl2I3w0uXP8Wq3peb6pylFvb0RjVu4AEUwr93Ut/hd6R
pzBzWsC2f+Sz2YkivSzPImPEHomY1hzureCa1PRqZdTrnHMFR42jfmxANUjXzJ8w
1uLbra4wHAZPMOA1JdgGQfNmmX3nayGN/2U1uW7jRn/YDHGcxEqpYWBQuOm6s3w6
8eBevqn6vMeSuFoZ1lAswHU4qKUrui71ZpjJ+MxkJVYT96JCa/2jqqNoDpzbXQi6
aAbrgyLd1L2OkbtVAG7rDsuyboBgsY28GGOeo8DWZkg4Fnp9gQVrBNih+DlDoyZk
YClT4P3ZXWmKwiREEI646d9rTugd8cujMIkoymt1beIpoRP16aag3gLE33gyk3hS
/KU1RoBQtASwcSMKwSVgX4HqLxQqBdxmVQ4zjPmGg9ziYQE0MvVSXTKrDG1fnIgp
jF0GHXAfyK/KpLqHJ3lysD3MALeVCLPuP0eA8tfxNcyLG3BcE5X/8NsnUdMarTT9
k5aNvtqWzz2ctZL3O3VDwiph5XTaUgLrY9AQHxZe1n2aW4J5gD/Zha++iVNTG19i
xcV/p9K9CFVUGZ3lk3MdmD0cMGNnkcuZKa4pSels00Ywo/gRzD052924nx80iyp7
uolC3QDm0Iyny9mFnKC50WovQMcse0yasPKAb9IrDHZQS//nPr7aV2ip5B2eNTnc
00GDEsIJ8baL+QRlv7aGboQzCCSGhvpwySPGSWLH55XGNMuGLK81ipHAKOCR9WTZ
OZA3tKWe3semaW4tebIk+Qc/IiLTMXeUlZ9KHc9Ud3MH0t64NUHKVfva2PM7LOE5
Y5sHHhfoivCoe01dNfSmNtRZdQLyUCPkkHFSpSKirekSZHV4cOoB4cEKRQhkaMwK
jambEKVWVw0AoOUc9PamOGgLjvA5elIgmWkQk0eW+bkPv6AfvFawhCbGrF/6Adoj
TOefWePbF5ZlCgIJTzFnMfMrnfJX9P3W1KqMiUMcQ9gISZ3+seRZAVuDmtikVckj
JhjXsRrbwfiohgyWqCbcBBQtzwy6YEg0SNHi1WDs9JybsawIJswZc6ePz/Rfterm
flKDuV4hnCwfYlF11Cq0i9VPURoqjHItEoPykHnwL41IPN++REE1526rcztBJ6ev
HMI1OovmkS1oNHs9mTbnSDJhgIBAzQLAskFKcMjPTqM8DceukxVf8UeVWMMhlNYB
kQWZfYAjGve1K6NeJhX76hUlGzdBKCcrR64LPM1YNm8snSfca5UZ9DD7+K59IZgQ
e9T4Y6lpGkUL9KWlMXV020uTRmf52a02802s0QOfAPiSKaGaVbbFafKS6h8n9+Ps
I4HIG++MC6k8I4WsK9maBWoYB89oSNf5s1KMvzbU0NIgMl8t5HV2HEPiRSKeLXpy
2Oaund5PMRDIC3+hSuDgivyoYjBuMvj9/tPLAwBci9thYoAArBhM1IUtDC+8vTLB
26JYkBLpnZoOcTtZ+F+0SjiO1t74vyEls/Rtey9AGr4X15CgUWRHGrM1CNwKLoGN
5O+ob/OePm1eCZe2cluYFuUswltppb9aVoSdsC3Q/u9RxayUfq7LG/xwJaXqxDwJ
cvIergHMobV+Xhts6mjVfb6fbEaLzWin9ZZC0AyqEQoTSlRqlMj7TNiJkog5M51Z
HvTp8lA3UnSeXWrTfEvBQjRD14H08MkF+gJkpYh/abH26KBeRK/lQF3F058o33nW
3e9eYDHmjJ41JwFlrFXzmDgZ/CTu8kyAKIa7Vc1B+05Dqu7IAXx7z+lBXQYCqFhs
taWqtTn2vOt3rkjwjL30LJaaUthsNSbLuyDoTLQwNuwGbZHok0nsQqyUGNZ5CRxf
R0Gfxyz5ZeSzDPkvf0cua+F2dwGlh9SoIOF8LzKZSDgnDl2w9TP13OCjdPYTdC0X
BC7Q0xynALfkzyr7zEFWfnfIs9XcGY5HCWlUWq00Gv/DNHrFNSDFtdXgLhGfj6BE
+6edOguvhMOcTO0sIVAVttLsWsUeHG750sWfI7aPBtYfji5BBKcPMsm5toQx25+o
Gt9MsdM0Ds3+HrXHkCA/b7l4f0DzdCvscM615JfGNyX53ZoPMhW0/woAuQwN4lj4
SSnY0RiD519hQQTu3P2Impp9tUHJ/8s535wG9qFjv5th4AIhlZ/IlYdsdWa7Txtq
pIY6+yx3jZaUSlfZPK+8Yu8Ny4Si+eenScpDIV/HFD7ohEpBmC4GP0VC8qEegmz8
Sd4gFFMuTg+Hfk26Hr/iP6z7UjuXu1FKE1+eCBLnRL9gUmbcCcM6L1OD3oB9ztkF
ETuUBdSmuCdsBcy3ZqjsviCiGk4izzfkhY6ihN5DZGidkLZTJ8zWdB4gs8dy1UKd
HHljLrUaQhgenZM6+r8Ee7ABOrgVUAO8CBnHdE4C08h49W+cjfSEjq49hHmIw+N8
NfVjzW4UoiUcLnz6yK3j/rw+DNyZ/sqsK2J5cjaPtN3tLvb0MNh59QiMO/pQEqiN
qLfN2ZqIgFF5WCDlLuD87uuhq0Tv1rlh+0WdDG9gCuYuOdE8CVGbsixDszgkWg2q
EIVxkStBs/giN5u7mP7pckqy+MBVLt3zLs8XnPlRWYAvhnHZpHERIfAXJ7FAqGRS
ZqPMEqZ1fnO9RyoX+eX9Z4E6P05mGFJLJDdVDZCSdIUhowXczAVGg7c0BSKzHWw9
QwtHJ4ggdZmTJLBsKI2L0yaMn3mHAo1YaE4tuNmg5Z9IcAGuT6GWRLO2COKdUioc
1ocqW8yAwxgulfzdJ2BXgO2U+k6F2bR1ZkC3M7mcISotNoIOSJgJOKkIzzPZluaD
FRnQIaNgrVdcN8P4GJ+MGJ/b6FkdS/C0FqFu0/iXonXJ+DHkniB/tOZeXbh58rab
O2WuGxrT9TNZUvOXBtEbiRsCYuRr1OrCcTpdVfVMwwy/ci3pZ09cOz5R2zhTiGFp
bwNU2vjhgf3OLN7bIX8cT4+aMAx+awJResfxAKCs4HGN4nKSH8lbHzX0pvqUi9JM
54VRRmKFT8Bo3o92s0zQfFfBuepXPvpl9dMqq9uTYvj6zxLRw6xz5IaOJ3CQqLJ9
q6YgForbpdDf4WfJiecKxC75YV48c85wEm3QtKbv/lfX7UKqA+ronrb8d6MQgn6V
rQPFq3ZRa+6Dc19Wsz3RrRha+G/oTX9nbOFLvWg1BapSQCUnAXpPQIxfMY+jUp9h
0vzomR/V1XeuOE/p4ZfHhsIR9oAPdi7D4pFxENI/KTqqlVV5/jMdQ+JIMpwHFan5
IlN1B8vCQsPqSZkjeHpxMp2V0NFbwzWiTqzSvvHSrCj4u+gSYXYrkIGuNXp/M2c3
Umc55k+Lfcg84Cc7BEj9g9nXnLjimuo4uSIYjhVD4qZohuPa/oUgfNHRbCudvNkt
QtaTrcaw8kknWe55Uyd9yrP5EmeMRyzA0b8LczjgoyLEUrsqaJgeSK3fkLtVv0p1
za+BciWb2gIuaxsbRT9dUtcit8/Y2MLkqHlJb+7UbwLFGm0VcWmp8hRGIQpKAWa7
AlMFRqmfcsIz05OFk+poV0EwW5We5OLiMVjfZUEh4mSAr/xGufPSLzZtjJ7JkpsX
4l3XC2uclnXogxHDm9N2gDZiYi/ZvUo3maN/2gUkc+RBKU8nTOsTNRfdssmZ4lZ/
FO7VU1OxzHFPRK6Fd0WLYhUPC1VbgXBHx5h4HpysLQalh6EO67WD1u3Dk2PwD5jG
fXkNpdZTV2x1mu37OxbA2jqrkrnUbuYZccdDIOtaBJR9YTobgTyNiCH/DMHfc7fq
JOx68QOOMvHABKcbNbzSelYmbWpNI8mFjC0l4wGg5HHXFFcNVjbOotDPQvvEvHZf
AF/tjMpLdAW1hyCQM2pj4gPUzrhAxEERKz1u0g7sekYCOZSaFZMUxqcKpt4HnJM7
RcKzuSBmEgCPE7auq5uKL6PH/PIysBfketJKAx9oHG57fFnXXP0W43QyonIfRpjc
MA5tMUsbPnGENEBOtzs7lIO3qIAnd9kW17u5svkUCoT4Zw3pMjWNxUtM5tZCL3BM
rzGjjz2Lp5KVZnLT1IxJrgJqwAeALJPKtlig5NBHeMA+OT8pkr1jGG/ZNbz65oAE
4Rs4pDtPrMomMc6Tqr9z/+mNinE7uEqjS+c6ivwNaSMdffufbIZF/3sGN8Kxq8NR
XkvZiBRFoQj1cZitqtMJLax+5hJ8064qWYZmKkFHNegBLgv1VRcnTvL27VA0uohW
LkJkz7Lf7zp6/tqDmeL56UqV2em/u0W734xvKUm2vQy7b/xBuplcTOZF8GgzR/PD
rSAW7u8hhhUufldCSqLsNrBL1cSsPAKBCkiscKZ6XHP8HIhF23Y/Q0jpR+KdKda4
guzfs3BTNCciZNDxJ8NJFwJ1+Mo5TONzEkkTmlnwtB+KAJJCalGboyR8KpWH41qc
l1vBrqH2W6I8y1GxkxiysBOyKc+JOh/em65NSleWPx06kIg8D3XpeAEl/GNp94ii
bUa+2OE6ZP24Jml9rOgS+hFjqb5UDUoCrnTyrze58gT3SNC/L2CtUa8+piN40Ywj
9+QoKFoQqWH2vbS+D14We5DmYL77EixtWCnnZxtLTP9SuLgLSAlMx4lOBuWuAJkf
9sDZaF0atToHDg5y8nPEgPQEozwmPfqumOXFGvCJe45hRmmiSmna7QLw9mED+sS4
r9fU8QEWRoyZJ7mZvxU1k6l6m1kEM8adYapTdh95/UzAPPw+C7Be0qU8y+2IGXVX
KDA/k28t/r55TVxKHlk/nXs7ywPGOvhI3sgZ0pokjdjeLtotOInbmF8URvvBpvqy
UeB9425IFSxj35wIzdV+2fN0GHOxxiY2jl9TEtbDfCfz3ExxNSHY4dTi750CWjYn
OeQ073s0pp3ud3rxokc6cbONgxXulzKYUyUEkk9lB/sAwRG9w3kG+0lcpF4xypbb
agbl1zQI/kQgBcQizqKztUJxY1LK4dgabVeDqM5IlcanzPqD9U9RssOcOQsj30qM
UPRBtVCZuWvzSvN1kppE1THn4p973OI62018W7EGHMh5qYEZRSlF6SKUQKUUZQIf
3BrEjmdUCDRsD7Vgp5Mp7gcPJhgH1zBM1GDyFyJe7NE8DtlViUTDqzedUFqInMGy
oGyToJZzM5FpdIqFwCr4kCFvqjoGcRp4gmB2/ZHYjG8NkkScz7MRgN4i/raptsy9
9oY4tArtuRK4y8otWYObQ48aQk2TWvQN0T6O15xjkmOlDXlLj42rHqD1J36cEWdw
PM6Z1XJalrWZHj52VPUpj3GcoCnPDmZzsv+Ti4daVi6DUkqJxIVS4tXllvN3eRpU
l0Rzj/Ts9P74msnJWfSuiMnc69Hu5+ebvNeBRaMY2iGFC5dhlZgiD1BOm9800iuN
WYrDbF9Mobhl5dpPw8TmmhThtd/IxrMu3MCieK/gScYkPUTq6Uy7sWH22HSl1EZn
jXBeFVLgxoTQNhOJNIvZs9rEQctzaoHG8b+E1EnfPFJtEvp5R2vmKG5L3Q45elT1
qrWmG78SMfeE9H5BzukO6YOjDAzsk1QfSrlD01HZoSY+CEmVg1BHVjnAiUjl1aCq
KuQxk5CKEuH15sUsj3one5nudQPX6fq2TLNLQNSgGAKVqvinAziKJpjch5u01CRA
TrcmVl0QMYafQ6eTDydFp+CEXXzF6brtJtS+Pc5lXsjPPMW/NGiRJ2dwkirlqRsP
r7MDtRyvHGVuM36IexKh1jBozwoF2IHjeoyAMFOXMXgX77vdTuhm54d5/+1KP7LX
yVKM8j3ctMurHGNSFmN99IBKuM5GIOT9FwkbgYb8Pm+oqB7DFvcRGsmr023fSVmT
zg1BvZVhRBSVuKrMAMvq9jW5+axXFYvJAc/GxRnkJQR6Q+R5HhMhojS4RrVameVR
w0MsHHiv1lWH0qwAExBNuIVu3XT9QfQKGrHmBdOVPnCyAe6ZeBzCCyQfXiVibK/D
SQGZos5UQpizi5uRb91DFUX3lCs1WPmIQdHP/tFJtWdQAt77JTWizNdLRY0LOlDQ
YhblgkqKaSc62WxHdnBE4dGqtVwZ6clqN+6PWfmPNBJrTbkUM3uYxICCI8YAFY1+
lu7pyoIxDKUyJ7nqrbfGMmnJYe5QCHaVrw+wWwsS8r0HPwwPbOXPVSgcBRoC80H7
s8cik21+lsXgCFmuFGoggTGPi9sLlep2z7H8t6Ek8ysO1qI5ee9M8w2M6CIJhzJm
YqfPDZ/Ty582xHutirIGhWdQor1z0dhcX06WSLu8r20/yxTnZ4YHTGM3OloycypI
Ge5xCKDtoLEc/07bdLz9f1qYD9+3dKUGKYJskSd4f0Hr41oi4qgSgeNRHAmXPIUd
GsFlEEAf+CiDvOFH94P1JE3IM9yfvAjDGyVMDRY0jqARQC1nFgLvVfVDrTzTZ1+w
VODBUCcD+3dURUq2/m0VTlcz/BLKYL3gBDf2Ugu8SeCXg+Hml4j72wPh6HAzwHnJ
0UDKEQpoGiBOYWpt+6N69II/2dCItHGBdyykXX/rF5dl9BKXkxHdQ0zVdD08UGo7
GiJvE9mQBYUqjlnTrKv5yqtPBZTNipnl0oaMEB4Tv4i51zPT5gf9vCeYKtTW0ndX
5WGqmsxNFOsqZy1oJ6z8CNYi8W+E2dm+HwyT3wK0dtMqVJn0H0A7kbUYmc258eOx
wOYdiD5PK++4hoS9HQWIdxiV+E22IOTtBVXE1QiRq82uq+DRlJDm0D7foDCIk/LJ
oLZjHxLy1Ih+XESkEaPRK6UBRQda/Y0XqY6UUhEZmtUzyB/JzqC0wfhxlP7I5eQf
Sz4h0zCDWGurkxQ3LMKHiKJcX+QYGV07X0WcurG2shX4+lyPeUnypMcTA36vt8kn
RXbzgmbh1cxbMtE4joEamyCZvyufNwgzXwZplzFboVzUerTj+za+ZvabVOZ3Dtnn
c9f7XlGLn+8Lc2KnWr72UBbGs0GqkehMzCfw6X1lEjaDqUwZz9R0sKIDqXA0LkZH
E+yZSy2FHiaf8uxpCN29jl69Hc2ZY/UinT8SFTzULvBcDBqE1qjuUeQey80syrOH
uWPripnrybuK/737hdBQBODkBpxWxD+oPKBuw5FHOcpGJMqOjr1blFoJ5j2JlRhG
VcJnEzClohEm6TxfSCCyGVB5k6G2pq4bz1fpwe9EFuDIHgzUfM0bybWkidWM8WXQ
Ht14mkxy6Cvhlpt4TJzpicFVaHz9KbzVRHUIZod86hbBIFLDrJIN/lA25vrZ1Ab3
vg5PCC42GTQWdPFF4XYmuMagdDj9nvfTdpuwL+qkmyvDNakA3D454umGbtHMhP4T
X+5Z32i90MXMD40ijblmiIrgfeEyDfhlfPG6OfQp89Reted06PunkoLoXAwQu5Vd
06ePY9hLT6xbk5jRQDo5NQcESuClD9HecQdEYdYPI6BSMP7FYehF3D+GYwWqI7EP
HGOqfKZqWLKVypj2km509Xu0Tzmn978VSZEuWLo6HvDMs5quKtM7NpnhinsMqcHF
ey2Oo4DghRHC3uqpP/Z4WJu2FIiXqpqfhTrHEl3E8GrkM+J3bVUBR3zKNXcvPABL
N9kFHPflotAZrmT512bPgJn31RNb2ML1cpibPeas1auw0n1HnkU2e1pSTcAbk6u/
p9XU5v8b4BysbfWrOplnGV1+NN8I5bRvGw1f6+tRv4oZSDxukdyHQUyZ9C+G5JDb
Wp3BKgUZTBoks432OQlefMXU9/a7XvWilthjoYaK5TkR3mZKZAfqYvBw5Qrb+lZ0
XB8Rn5glk/OsTd5H2jTQNbT39WfRzGnwieNxpuK5U8WvRmJs1KcWOOZijsjXZ36E
Wn9FM+jgJCBpFe2HZ5mGPyd/KoHjfdUl9k5jknI0OXzxB6DIRJqPAMUJn132jhSA
c2qO7nwR84HT5zEfv582FY8GOycFRVRoh03mYPHDF4eHMxmwkhrsy0LY4oK8Eb/1
7Q9Bl8aIcgEfelchceVlWazmVS20vePHAc1wyayarWbKo1etrMBQ0MplGprkNc39
aI6HRcgsB+nQrtTEAR+F5/f7xY+FC+5HV+5Qh43/kAq+OvCqFbTPM32s4Te4w8Gc
TJ4mTNraiNCjWCaB1nDZqAO+sjx3/hWQmHitGlqczbGRZ1p85Yt49DcUdRTaYSVW
xuViXIdxYYyxShhmIytjs83R9px7j1JtYvQuoyYFF6cNNSsTu8icG22A4bj1XfVz
TH/tXf7ynNvXjau7poJzZVubLonQGmzOHyuZip2lZJUDKY4czzkS/QmOFw/HTASj
ojzJwvwxdqxk14pZ7/EyKlHdRSsjwgfyXKC11w54RR3XLnunOpXYmi8EdsrXhKRF
qacwa3ZzAUyQatuZBzVMyapAs9+3rQAdyCjfRoz+UedQeKVIJqYf8sdaETiEMk7l
F/25DtQmbQSkr0VMkyDBC+JyXMHXAB0RrInzHHCs8TV6Fc9cK5eh8Or7CM9f0RBG
bf7xVfz1A3TW3Sou3NVrKQAc/lI/Qrec5ScCjOo5IP+iC4MQ9yS4ZxokUD+TduMD
OA9DJJoNtgC+ayqA+cw1F7L4nrGShhHtJ1TUXUogspyxSxN5SgD19biUe6sn7r4P
TKLxUTjqnPExzBw11S+lJKFN+mLSwX7IwvBvNp8NAK4THEZ4hoT9z2C1P+wWmJNW
Fea5O1f4qd80nQjS7EMDTT9X7YgZeSrYCCRyahSkQ1sBTtm/sbEJHcbCd1dpI6bW
lV5dJEcIaRGgbE1O+aSMbkvRs6ZgrALfutCaZQdbWYTwM7TmjtOtc0nYz+FaRzQO
qxrOPg61aPpx/CMmIR5g2sTnkmmuRJi1Qr+bPTBv75jWFkL0arGPadhOE9IG6XfR
SRP8c0FZJDbm4fdbebB6Q4hEITMSXA/pDRgalS2LkK8VwJy2W8uKsNwztnKTKzXT
fguzAHoMcW2XTPdfu+ctoUpMi0nlwXhoxtKlqSUIEd7an/KXDBXn7xhdrot3uCs7
d96SmHB5cRdw8EfbB2qB4YUU4kWvcEyUhazVT3us06bMKVd7HfoHsitwZfZPPSZn
OHjl/FvQWXtb1zfODmQFjF/Xcx7LsZrDrcq262Z4oIqi5hRPmXTyhRCyb4tTgEqt
cSiCXcFp7nBXq+7jnLXf1i57egaUPiII2K7S1XYzOXc39L2p2Oc6ZZM2JI2xD8qX
gbGvqxSW8QmLm6Jf4e+j3JLPkCDg7fVpk25vWC2dzaNZogkH+JtcbXlJ79ufBAFn
NdmpoC/5RGN6z+IQhc0c2fTCjzprrXQKAfk0sZirkHLjeqhS8B6mtzZh0JTWmpBK
JrwupZQD1Au1LRKSdI5lFKciAKYAGknkX5jp6aFjVNlPdYybA/hlzN0M930b6oOI
fVBlgo+ir0b6ky/dj0azsZ0idqOHrOx2rWUcOKzl1MjKBhWTMgpPI08mnFJTKwyZ
+RGwlk0mWDKd8fEyW4lHs5DJEzjW8Ojo2uz68Aax36NaHfIneFJF6T5J6QXd0jSF
a+4FW4keGXoVjGhk9ed2px1exMwn8b3HDzmbYBrJaV/a3IKy1wzeXPOXrbX1IzVP
YWeLl005VPitMtIl0ZLITrQLx620yPjJkH7qQ/of5tD0gEOfTi5fP4mjrT2oHwrZ
3nIV99flmBuwvVD6DWWg7cTYlveoxOCHpwasPBEV2zGnyqwH3N87h/C44qYK6k2S
pKCujMH2zPTMq7C0rAXUpQMmPnS6degDyKRltS1D92GJYhblw+vDDkAEOAt7yXMT
4MV+lPaYrpe8E+9LUx4kVK6Kz6VNkmcY8On7kOd5xueo6CiolLlycQjo/eYpJh9P
i2iNCwvXYf2z0GPmkCQQTRyJiYUb3htAmQ2hKxV945MFhoemdJdDxJXbGCJtPfTi
mAGBn6rpu2Ivwvhtfo4o9fJ6nrApMtcHETcYKiBAk9MAkktn/7X1wZ1KmQhZsRki
aWcx/Z5fO1jw69OxE9bsaAUZqzp1vt38+tQtCZVxynnzmni7P+8Zun0SZLPSBl6t
JSRiEqB+QovkgEHalVWIXFC2JPySGDQMRZGKhvetdJxkci+B4I6AeGUfiAxqPQbt
u3p55lxRZlnUa5nZDPTgRhTz9OYrT1eod20lmhE4GywUWnbfY6N7+fcPzrRn/g5M
AEg92IDQugHC/Om0r7jEvhtJf9LWJuu1AU3rHnSo0WOdYzHi6FK8Cv5MJ6z5GB0w
OR497KfA63/z05VQiKZcgOKbhTIsW/aITROEUMcTkrZofM9dXZ0FZIPUdLd4lvdy
7KyLwGMZHL4+oEuNPsewCG9ogqpuSQr3vrwkwPdHTlCsA+dIDv7ciQymdFpVzxWz
k/5zQyaRSaSxlAhA4gZ7v7VDb0e7uafIaMlEAqgxXsnfKcrSBuaEPA8QLzMK5bIu
QaopFAZWAuasD0UNbNKHwAWYPSIEmJwmVuArbv5umCiGPC3CWCxZZ1F33VTtQXu2
DrYYzh0zehbaxP1sw8YXdix/dMo+VMNLN6w/jaw+v/SXE1yoVC8Jy4oNnTqerV/e
n2OsyTM7etpf1PwJDIg78qlI5VanZd8iMkaEHVnvaCHI54rqatI73/3bSpptyEgR
mRkyeQgfFqYnX6/ptyqY0unLZoT1Xa5hrO4fZeOc/weKkHusA0/4uErlrGvFU5F7
OHCqz8fyAcuFfFJziFQYv2m/pgpIJbMuy+khA03hl7VxyjhCX21WbKAXbsoBTDNZ
4j7n6LUIzdojFeKYXm39gO3BeYvXDMoll9KFNYJWx+StgWFgVnqqgiceYQoB/Jbh
G43LTIkC+xa37Q1QTux9d59pNt5QPETu85ectJOeOsKVM6N14rzggLvtiOS5ebaL
gu0YoF0t24DRdlqjEYfFpec6g7V2EDqQJ4IRIyKCDAGA7tTBhy655jYPs1SoD304
GBWEHN6nz9dmzxjoTxg+v0lQ8mhZOHmHDAqF/kCSjklNEw0m5AJvDJrp13GK1Z9y
nzbTnOSmckoSvLuEgodW1YafeUw8HjiRD6dR4LinDfY2XluY2bnAeo13y70J0nTI
6Us44D2BLcgxo1IvibjgZCoR1sGszJjNL3YTZ5c5ydQtFGeDFDTT+Ym8BoOHWY5u
Txnv6/uGXQLFN/rAprt2SS4jI72NdgLrKastlxqaWHG4i3ubR8RxcbCk0UXLWgUk
6a4c1I4NBqY7LXzUWtCvZ9QqOPDolYxd2j0hCwFqZl+ZuePjRSatHHWMlL0MFECD
vbS1B2U9sPkfXRnHTyEpU/0KXe3Fki0MygQ2fNU3qP46eYNxdRcDtU3ZrpLvqXat
bSIlP2Nz1eEK2BAGJxPKw0IXtcmyrLunWxhWYbpJ5UMJwOumcMcqxqF+/iy01LFp
l3Rv9gohlqdQUXzXwyFLBYP/GHmkqIN2wBMNYEf0LjNbd8p/SjhQpvfzGYUJ9mvE
5Xc3lxEJpmHKTouycqvnD/iunQD/CSnMTs4UsuqXvHEtkeJbgqU6m5IOzBnyE6Sl
EMN8s2/NCwJv/72QiH33nkhBZrF2z0v4YLFBD348cELARSG/X9Oll5x8TaBzc022
m5O0bLwnh3p5RC803tPuugaoHxsHJtdeojcyyqTKxUAfwdvHjHblFpuROfphDP5t
uFnWdpWDLOrAldtPQf+kSQ2GfzbKLzto46xCve6xS0W9+8SNveagXsQ1Mf4LHcwB
UmDKHnelsFBtut+RdKZamRNW1NshIIOYgfxn0F/+ZRcdYN7L6gdZfEpPZzbmz2Qr
FOvSa20cXjchZxNJGlOdsgZaIQKsPMH08KYs+7Vs7Kf3DQlnhnJ5AlEgnarrpECf
lQw94c5YtPu4UDGyaX/qxUk0Ssg4WFKTrZAhFcun1FtMjRf9npjBD5z1+ee6aI3t
BVt13QWk6OU/859c97dF91TnvhJyzlXA4j74ZEj8hNL8QeMqsNM+on6csFo9pCyv
dhoENRG7IIhrKEBsMg5R6IxGiqYeEn+v2taV159go0kOI1USTBTuvheoJiMT1Ol8
erCNqsdmAlD/GyEfrUBI+Wow5eaGGJGez8xsZUvFU9MnptMBR2eRzHjpxVg6ylA/
tV9gxR80gA0tzg0omST3J2BMTEUPFQhuNcs96VrJWM4yDX/6anuAqegJzg7S2M26
mQTC+gBoeXMeeTWYHM47ME2+Wa9BzAB99LFHTWRCX7tgzlTSIEArwHkoXl6xsxQ6
FZ3vre/Z/ZiohTeRuzdjNPMLqx2gW0aK6UsDBSOlbppzXs3SXpfAiRRv3XVLOwHj
xvDYs/JpcD13ZnrdVcp6aUQ46kLGGUj7DOEe3dgs7ZTElvOo2Y9tEHdDDU5aC+vz
zBF9qEf/qLZtD+7/kgLBNYt9pP9bh5ROCI5jZ5+L3MMzTUFEGZQ0Rd1sXkWyq1E/
DCSdD0mZ+Kp+YDhKi8HOFwmq3FaY+y70zh54nc/Ao+4b2cLBSEbg5ykLaU9vlv3o
vazp9tj1PZtNetCgPsUtWaqe1fs+u9KjyKR47IDIWA5VKzZ8u+Sr+lXZJnsvWgxu
8Wn+N5VAMKTU8ukHYqSQtvK7RfE6Hb2yQaF2AunPrTuOqtyQRQNpPyqEhfiPGsEM
EWD8KPGr+MLVtWlXdqTQnRqIe33323ZHeqD+gKFnIlias4tF/B4uD5RikWFhBKzc
nCqy6+l8DXVs5Jo/zH0JPQPU47td728guO689XxHzwzQFZeKKpSWTSvu9KspTJU2
1yKhzTln69wnB/plCvDOv/3+VBCYKVIxzSwfiKLPM+gvsGDtC/T7vkW3NwyTxPsS
xjr1ForhYqMYS5KPeAsXd4iIsiofAwVhuf9m7sfYKtrd8gmsbbWQyfS9ESCd7axj
DZzLVKu2pIfclYNESoAzirqFgVzfEh/RRoXzUmBbcg+S4Sto+qZrL4X1NOu1UaZB
XUiyKYARag67oj+TXJxjVgwxoHKqsHFrZKvyNVIr21RApvp0Hx5mJ9jf93E15JdA
I2TG3SFAOv6VsWLxyIKb00hvphQbPNW5k7zMMm6zql7EIw2xGA9v9laeu3JFwRFW
TO/M642yGnORRK4h5WT+h5ol3Yo42v3iC99HDz1qKdWr2ULGv8u0aBhWbOLTdR7B
N7JvPm/7PpheoTyJqWwZt49M0Fic+QUxgvc5PjU1qUYoWFBXkSW7QeKrVit4bb1o
bkGRER9fBp4faadgNx4VekG+ozSGpfqbNVlRyFS3heJBw8tG00kUq0ATIjOclnh9
wvED13iTd3XlyQStYbIxlWE2m5E596OPwxngWcjGM4h4i6V2mn93VjhgaRLpdtTc
2g41sf4WoywAlbCxbeg9YmvygEYyQhVJeMmXRER59lyyYkAmjWfOkSNRo0lrjGPu
fcuhR5bgDDRyy45qikvmKSW5ibw0ZVljyUqawj6DRwP1C4fAVFLW9H2ZXIBYAPM5
KjVbTO3dYuRB6SXRQ0Cfwt7U9jhBCQbKgBLv+R84+LkUnCEhEYeiSJRaQbjfWTjX
3ztjv7ARRHiHp4NKcR/6X5cmnal3UmrnyTCsHgXvfPy6EgpV6f7ZILORB3YP+GhB
MxbB7ikIeARBxuSQDVwwhdxDLxchNfqqWcabxqNS4lyzCvd0K4E5zMsCmxxCchV0
N9Md8U/iEIoM5G2WE27T+5aD6EfThw12Z0flLrBhJzPTxrSXm2q7iU/0krv8DRjL
hcFexjPoMvbHH16eKX4loc9PCS0vtC7EqfBDg2zwHZSEntlSoAY9kahLBiTE8GtR
uITNdbusCHXWXOFxcjU2vS1sVZw26XV7w6mP+reGjx/w4FZWiW/eaole+u8EzLyh
5zaGrxCq2s2O8CaZ5hTv1H0G3RtPX9vk5Qam/6I5EbftmmOrhAUENAb+cez1GUHi
IuBaNf1zGsWBEPqQ0z7mvorAq8q1AyCtOzKCqIW7zZZiMM2lKBaFTKsRzVoWDKwJ
l4Oe9H0sS7F4Q9VRr4EzaPAQL3TR2z/R60eTUgpX9xHCPlZPkHvne4F5OBIOcJtq
dVYuxXjd9odKVbXZMyWQ5fssb6PFVeS+939uUPpxJUMFK0trUNH+90Rn71Fmyuo7
T2JM0OgcD+N9Eh6QCDtXjjrJEy39Kgt0QyI6j8+upKmjdbtBKZNL/xQlpirVpUgI
Ar17tJf9Fot9oqfnm+CbanedQ5OKS8mQDbzfWYsY6RfgWAxhz9mt1oek+PoSTXri
YwZQTDIMM+isj3fup754RY6JiiZxtXhpfgpnSv86Wzjm3ByZJG+MEDI5PVwvHmYs
RTGrA12dfI09FIY9Ilxx8u3fsBA2KhNjqitZyOg8f8isD4tAW2nLJn8BdXc8nopC
GWWoVWEO/x9qPorwWrN0mj6P0PELQgm6bwAGAtvJeye2LFvtP96wjewq820Tvmje
ENA997if4w7t5EtnFqhVwz5C3WcqbN+M3ZC0v7t5kxzWODcP/R+qzDPyVzrSi6iY
a11SnuVV276CC0OzNqwAGpoyLEBRHf1rSTTE72OCZdb3AQrWD6U8UXdmDujLfne6
Z/p/0a1l64iSbS6s14NMWi7NfNEEZZfTmDrY/TszSDsnrSwulHkqofW49cd+lK8X
pNfbhoEukuA4H7fTwR/xZ6PvSOSIh9aStAE2OcBiraUQdcKSLUqMfjS7/af1qJGy
cWWakgVhFtzX951ORAOyuKShZdKhtZ+wmJBFq7X59W9RtBjL60KjrSjQCFbkDvFL
FqifBw/7RJFelAiFOcJARpkCws1xtfiIG8NQ3QzPTO6fDOeyLt2430t2WH2aj4cX
YggDlhCkXzArgiG/H2NN0Z8lwVbWxWau++w9eNHiB+B9b33HI3tSN7cnniNxCQki
4iX2yJdHak2DamCpY62gbxP6QA7OBgz31taSLN2XAcD1dmoVsneldmvyBbnO4BH4
2lIjnVRQs1WjLtEe8hXxSnkp7ixmPOqGv7ull7hb4ug1MTwTUBHnMQ3r9/cpPvYr
0InrhfB31Eztq1KDCmXOD2yBWEDwVANmNTrvL3lXuN55IIqSXCszUziOgYrntURT
M9U9Y7fBUGwLPS3dyHAa8nG4Ej5b3vs8cTKkaXTmy47LuFeDms6uII6kNKzPD3nh
btKtZEN4AF2RqJjxVg4gNLbzujqGCecwaThb9x9hlM1saEgPYHUZMoRYsCrclEmp
EViZzn8vvPbqsoyWP5yx1VkLu3T460dh4byUnsQOEmqaAFNmmdXuzLtwblqEm09l
DStp7wGZvrXoseFvBSyhVM9Dhsc9hxVJH3wWV/VQ6UQhTLs5fN2u/cSvGeLnvrG9
00mwviEHRG27bNHOX9vhqlmKr1Rf20kKYU0hXzahmFCPKFgQ3DFVaKl5/vO7APiU
+bxZVIA6JFjkc0WKCdyaY3GGL6XCDJMLqQJddom1f0LU6rMzmtTRlMyvZDQMi1JQ
Tr1YA8aS85d3KLlDRh7i6s8P30dOMen/edMZ4S+8Sc/QL8ETGY765bVk2jHxp6bu
1383Ez85Obhq56U5JumIevyL4UXi8bC2BS46Y+XRrtuQ1zFwBfq7CRwsOiY179Gk
cdHFazb43Zb05NvTkQY4HY43uLs2BkQMeDgt1OfWIZk/vAjIqy3yUuq4Vneqy941
7B1tkPysM5SNWrN/l3L1cE8M4hKhOXVlGthTvaukHzUzLdrULx6t/z9Id7XGlr5F
Ft1svS8Xoyg8vJiyDHvutyYBFogjZwN+wLe+w9LlyYK6tPAfBqB30Ii2mbzdDTpA
Q98Bprndo2dEoZg1d3C0mtrs23Y/3jXChdco4broyhjzwtLLIwB6h3rKjBQk6YzR
Q0cMKt5FXetYFmvuJCcfU75ZadlA2VHp3e0m3ClNQgMBgd3+b6NP0d3se0bL2gx7
mV+bLsOELHaAmX07s0nZNzlF/xH/nd5HMWyOdHNJ9wMERZ16MfV9Ck1RqLAKLPcH
i5SpQ+LBvzBEpntKjlfNdjqyreeu0CoO1EqjLNQRpvOEqEy+F04HWmXotKigpsJu
kxc4AnzleBm2AxL7S9Ci4HcflRJtqXITR6hAaWv9lcSl7Y4gXFnXJkKDN5urxhTg
bk2bgDsNC0GDJeKHuxqt/ybrCw5zdlzuKNQT6NvyjyA9Lyl9xIFXWEoM+1wX11ve
4tyalbUb7nPfm/nRbKAKeVx7PsaBmGDN75ILFr6uDq8KjD7t/+Kox14BzfWQo7PX
c1cE3kN8yozYROn26389yum+i+myFdcKgRUcEZcE8y7NopxpY2VQy7FqZ9icLOyz
DNOtnUdxu6WyOqDtjTiNVYc8COyAd/ibiCz0/5VhiFgzNVFA+wLSYzfC2/+Nukx8
pFj7uJWpZufOjvPzQxGfdPfV/EoXAdREoUri6wgy2AbGmGVc7jmfb83GJFZFBYas
57uAWUM4JnIvKyxnwtpBrO56D86DgAL0mendlvzA1pJWuS1FVUTbntEZqIj0+uFt
skfcRtdsRaFtp5uGM0rLQGKzKUl3/KrN9LEDgfrxli3eEA6D56hiKYneU5picF1M
LGt9Fi138uugNVYCRPQIox6t0r2WoYBgMol7q4kCx5JVhI5+vOLoG4XCOSL38EJz
zivy2pHtC3cYRxnCCmSkU6FTtMEFTQ1QInIljqK7vJgkq5aJWbzE9XwPog6ybZ8A
nxjV2uHCLM15LQQkRBjTStc5wHwkP3Wkggn808lVNbRyOGOadXzpHI0u1av3wQ60
Zvuw52zq/YK2emL6hhGtvtguy3LKun4m4XUqyEFB9NQ105Q8xbhTXD225fMhubbi
A+9rNgguO5P52Tb8TIeFjjJRzTn6m/GxqCupU2BAKx2G5btCP+4J2PZlX4zA/Vze
Rur4UZnw2SPhjEHyP8NmzH3YIGlCxrRhyda5y2+uY7RuKg/V4VnqnRMyQZMEsIe1
wtPlqYyCrUcpRjoO8hAC4dPqagA7A0p74+Jv50eS7Y04mAa0n0xUpchoku2xEur2
0IOTNiP37f0ZszYZfyAYUXl9LuAo8S6xMJI2CyTYS4dVNYmwatUnTqz5gWbbNgS1
cogHx1qrjsDzQKrbyIQkRlpmuSn8awyy5v3BS6Gy0zk/opZIc04SDMWp/mRewq/r
W8c9J6teLQN/6ZcI/w9VhkgkFNFdnhaHCRFGWjUtlfDJBzXj1Sw4F9UTYwuj56E9
5z6uPOV2+qZ6jPwm0Z4hXNbeas/L9z1A2s2GJ4fMg3Xw06vFImUOGCnrsDP+IdrY
IHD2KeiI7oXZFhiBsGjsE2t0VltM5As/i3gTWHRAxB/06SK2qSSAFxiwJcLbh3OE
uduiMyf9/xJy1SIJglA6jFmAyK0BGigjAced/KdCMgwU7QDDz9PaUvDRdhY5etvw
9Nk8zb6eXtkoa86g21r8qKelWfTKqwWgchjA0nzwlLXAz+7wBjLJ8JayjEyGVv/d
STymIf0dYFwiEKGsIUg0dHhVoK8xvlrchsEtCdwbHCVa2z1uNoC32zIISMGInkUt
Pnbks5x2xPzOptU09LuJNIQXrclCMdIwwy//z5v4hvOzyYZ/8vEOfbv6fRHKrLfi
4q1FyBe7DkrJy8IUXFEffdbjPAPT8tXFzRNzBCmTsxUJsgiMyTFSxG0kLu/7/kER
yHmar2bIJnOgQEmT1Us2JdvvSd/a6+Bspxu7q/YBas/ITSXSQOi3QjxcsU5iUcFv
3N+CtLU5iCjwN3hXUwuHBJABpN+vjxBjyKxLCK3cmLgYo76HASlYgxOAT2hLMbN0
GlBCf78msqCSDOxzzcQf4OZ13aS1f+gUOAJT3LoLzKUmzn0MWR0QGqSf8O/oCPqV
SXwwmEhGimHAj+fVZupJlUgxDx67Gk+kOqAe54Roxa2lGza8numy1FMoxa3J71Uv
7BFP+EVG8UayA/MyCtx2rWKdqJx2vLYVfrc50y2sxdPIY5ItfhMxVK3nm/4+tCF7
RPV4R5bvO38mIGIWsBMkvxR72hoMgDHPSGduwFkHnIZ8Pr6bAHjaUZKRZ7t9L86D
mGjIkp0gM5eq0ai4JqbRK0TYZs4Hzb215qBMHhl2cg7vQcZ14kazNQpd5NopT4yX
YS5sbEd5ri3nxVeBhlwvy7URKD8IdSKkx+fmFWXQOtCLTGcUnYLrM32KN/jm1aTU
bwKqO6fAVw1XxO1Q8aU7woi89fMd89ihmp8doRT8i01BUCWqT4XtP4U/R4PVFY9+
Ut8T29pJwyQbv9b/VaVGLhSh4yGjvQ3yPzt2VU578S4P8NBIhbz8fatJteK2j0Ns
QIGG6Fzz9pzokaS0maH7jT/1uWjBgH4h2PXxsmk4HEXYGXwO9d4WhSgmLkUjk/95
jyYSLiyadKsggT6oMJqsYIywlITxv4hkOJVpeDIeek/KPAMxispjILguVtFK1bsg
WS3SQF/Hd3d267IeVRMoHYDfKW6Rh/nGh+Tz+tn029ppKYj5dAxfk3161m3PmiNx
mvVIQ3yfmsdXW0+ew8yGyDtQLFedTPLX/moz23B8L34dRQo4aRL11hWLPnWFyl8r
eCXWSYZ0J3a7x1eCtlSSxF7x1wVigehdePcOZ3vIRfDeA4NvPaG1ngNf0QfyMThQ
pNhyoBZSCVGIgr7yb7VSNetUNHgCyUneL8g2BaU/HckpCDcXmAQYLym3PV853jIM
EJG3f0vBp0rVz01+IM4NjklYwNmUQr34ar67Xia9dupWg4e1O51BqpVSdDqoLlg1
Z790PWx7oQnMKAvyYiLe8KGHruJHD991E7Bu5ulHj0zUxdpR4X9gaqlb0f7prO8K
vJwRmd+19oElUlOLo3Jx8cdsAYzQGgWBpAaVdNsUfvcshd5lrTkOdiGRD/EMzo07
P++eC/s0Il7/XnY2rtU9/m73sFpq2vvPqUrm2cnnM0qns4NUREF8WOHiES/6qCCz
d//MBUJhAVRU8BMdFZW0T7QcakkXBa3Q981C7UlwCcSRqQPlCU7ieYbJLhjP1wFx
2ueIaZ7+XBEuoN8MymakxZ6is13ssfxQ3losfI/LcFa+iJjdGj4Iriy+P1i3CF7t
I3xXj+A/lj7Y+EIjea+RlJk4RKtUWesKXGlhQjrsOBsp5Bt78QtzptDTp0rBpU/i
WqMH0tpzvW77R/HqLvO+qP25UMo0eGhQ612HP4HQFj0dzfNDSOOfUQQbm4iM85n2
zpr561lDz0eDu5CGNgfC8SxRR4xChRALLwkAXtKZ+99QC22YYDGfCZZQh4RQI9ps
6uk/An5lAGc2PGMR6KIIvi3hlB99kBi/YdqxZHYl9sslBAEQleKtL2bpHHSl8Sxp
vE20fyvJezxy3U2kRguGRw6/0/WrnnkHkmkVf1ZmBEEkhbKznayD7DvEZmBForOn
femYaiYG86ITTp62Ivp/mzbzEqpp7iD/GImE89eHRQXjDpIz8CeCX7cyLF/c3yhW
GjoN3LYy1Y2PnqL9prcx8liDj4qbj+rw6R47yhs18F2gRypoiO2tMbSw/i+SIZMq
X6H3nFHztzxZHzxnSVKaDeZnWpzs8/uhv10FFjcVngEiuKKi/UbReHsgA4Q1wY08
UlYl5J5A0vcSvcdard2GD8H1gO0HXnzMQRdcDkozJdDk3YaYRBtvL7hXCpgbQW6N
Sw072BBFqqy8+XXDO1SLaMDPT9/zpPUQaPAIh8IlPakggqWN8BK4RnMgtzN+litd
iQtHw86GGE9274d6mBwle9MXODNxrYYebBoWlC5KF7tbNz8Pkzqw2O5uf3V58efT
woM0b0dUMTMefhrkRdv0usZOnyz1ulhn5R+qWQBoIAEu30n7dPjK3I/m9FBzy9r3
KXjyydMeZk1pxmTpSiEjwnbG/IAAoX+cZAt7R+iPJKUZ0QqviB0A1gf4vtnwYUed
90gv5Nc5y1C9DIotCUwBc5UEghYg2BSPUsE7z1sM39EREyFo0Bsv9X3/MzMmG/II
YgXCTwShNLEkALEwZe+3jvva4pEn3/XPEWlkIVhIOhJm6RuFnhgKfPZcXF2O8Ar2
Rxo10YZxE0k9lanWpynVaPBfgmhcDv9Z06ZyS9zWEKq8fztgdooH9wq3y/r0xlf+
4AQIWcyatad7lu1kdakZPf/LOoVqisfVuiEe3+Rv7bFi3O4hnPc4/ZGEbm39FYjQ
V8UICW7WtfYODD8unKNgxB26vGmZstXI+zO1x2AO1SRCQ2WfpJnQWD5pH3w2c7cq
+Poa+dFcc+pRoaPZKxDreU5N00i14TUMYAtmpfMQ7ANqBskWa92UqyaKgqcsIo5f
wsThHZ0Jz9Kt8CJHTzmAVRondTQQ0PO3SOH4zwZXSvAcXvCQurLy6TzrfqC8uqJS
A3TZi9vdXUrFtxBJK0qkkZc0HU4nPLBuG1dk7uecNUYWoY/YZqI1Fpcw4Yn7XMKA
SAy6aYZRyPwgOzRrYilYHB7sosUnK84CTek270DW057N71/1sugZJilzoIiTQoZX
xTeHDuxjJ9/XxoYZiUyFm9u1fVNv2v8KZaZ9l+HcWvMoa6Kc5lb13NOmoW5ElD0N
UHZD0sq215R8Ybry39LCnOstKQs02Lq5qOSHVXb6ivo69t2QIG62ROxPA3t2iyp3
dx54MbSziwqAfj6uTaQZgz8OiaIiYfweH1QZKsntVKqHn+olciLlZR/BnIYRGRAD
3HOxRoHuzatmiNBb+JNXbwCeE+Qzv8ibmKiYFQnIRsUvk2IIPRMT+2ZdfFEGgaf3
WB+EwVW76uG4ecffAV+5ZmFzflVCoOlGrGzZz7TQOoDBCSrb5eonVluL9VEWh1jO
9jT6wcdiNkJ6Oa2PhS96a1ynijfHOzgn2+P4sTMuQQKpcxGaXCmYsM31XMCr0YGJ
uo2XW4C9doUA5T8o0+WQaAAwqiHe8fhjwmZQNdfSlP5O038WhyMBiNxCNID0p+09
9jpFJX/9y74EZ78U1frfiqLzNVHJllZ7wGkePDl1rFjtohYt/NoVCHu/LSBkJYE3
wKLYHW79AvtWJV2e/HvLiSvXnZComb4YDZgqn7xONfzp1A5GVG6M7Pcj3lzqCgIc
dXugevFDA+R0cf1RCQhGuob+ZMl3X2Al2LzfOUQxv9EMGhBRQOqCoSayUjXFvlhC
2H2bCxnyO6RPH4t8cZtXiFJnst2KqThd6HqMhZQufIU+4t5hk5B/dX6A0RrrgRma
B5Ez9GxqVzdfNOnnI225rvS0lqtseUXhG9yCeaP3uUPyrJlL2x9jvbVjdaj0TRj0
qLd/0/IrYubDxZc9QUm+PIcz0xxu72FA5jtin4MGoLE6jwvQfO703ZCgoGwgn6oE
f6Ni9YHgBHCtLTOp2KSxpegmltaCovYPUCniDhXghn9xfAZZX3hLuBNYcS2Q1hqO
zw7r4aEYwnbcbDrG/RVqmzjsWYE2Wzj3yJ+XMDmAWKXMz1W1Xmwbesu3xsaS6vst
n1bQ6vHhz24iMiUpq49TDzjNyICB0fbvdUMvIXNaRiSm1HeoIDFv4Jbl6sYY4KYL
aV2WwZW0SqSoqTkjIRsxKhkg7rWDs54awZ34SCFgWrpYKb33MEnGX/rCEyroIqtI
s5nH1kDrPeh5jwUlZegSWjxUEthaiRtASOL9wXFOOldGIOdsjpCwD40JvXzz9oYu
gNMokd8NBDZMUsgQp+EgM1zpUW1jXqKfNX4+XhVfnrWMQ22UBMY8KIxJJlLINaoL
3sBrqxpsjL7pNsvDTRauWsCoe0FJEo0y5nHmCgciK/wl2u8XgVvbvJnU5u1QWFmW
DvdQhtOKDSt6f9jBuzJJqSiM3YEKgbv2z7wAm/XtXASH/tXLU0LWkgj5CaYI4Z33
G0lLobWDGgFJJDwhUVE7qq6g/mXAaIo9ikZ+rO+L5jZWI1EiWPKbZhPL7fCAsFXe
rWU74ao2diHq4CjssRmgz0D6Z5mCbCU8RRQtSrKJzwROhmW2iElLWzbsYLeY8Cls
bcjwuzyCQFC5YS7AODhaolvZzPzgYOhtal5E4RqPvyMNblWmDAj9rmEaunA0Ex2j
edHVEFrW3A3ElkVQZ8UUL3anXDlDdBswzELj0WniChaZL1KzRK6XdUKPzU5z/f30
LW56Z8cVnGICKX8CbkGYLqRArqvk17AAI+FQg61NnVy3X7D9wUVkE3Gj/YHVZqZn
Exqgwc6V3AnEst95/na87VSJrWR3sDsf4vYM32hT6eKjG0DN6dI33iG7JBN0LGmy
KB7LZL22gGIEcaYFAb/qX0aEAHXd912WnWdvlt1/7eXqvaeMFboV8IMySYdJyDCW
5/Wa2s7vGKM4Quh/iYLEMTVhg4jTncMsUJOwlv68As7CzEpZTCTMM/hZUQWdRTok
wbpvCrEIOz2h93H3DN9xyMzsUg4hXI1LDHIFiD9oirxITN/kPYuEkdqPB/il4IQO
Lioj3G35OpjYc8G5DuWN384I+uR80emmfSHZdofi9eoDubhnS2C6zT7IkcqCgbFX
TOzmuZR0mbIa0iOF90Sc6gVVHQd/1W9r/2p0r7laB3b9uN9r08mmL9LmSjc72frl
Nj6Ad7wB0YlTqL9+0C8kfkCG1rDvKcWVz1+VCRjLqLjo1lRBlu7q1sRkopZ7iURY
x7QmYUUpObt8ChFsqcpH2sccVBeFH7Wf56hVXWdJJM+WecmD+WN8DtpmTqjKEjKh
uSnVy/gijsKK8uU1VGv8DEabG7lgDhs1gHcct6NtsFja0tqI6grVs8+YAuxsR527
5ipxUoMJ0TymIhYYuy+l+vPna3zpLIj1SeBWX0yKp8mbCK2Q3e/JRdpTooohOHI3
b8tb/0cO/+YsVWxOya7rP6reCIIjwEH7O+GrKBjso+v6bSYs/jxF4R5ZHMq/pszF
9tcYEH7HT2oi5cwciiIZ9mVSlFkQDFZmLHX8jVzoWVveEhaHg9vPptUsy0r7axq3
8gFbg+uMJVSrGIgdPK0+pVc8pxHQk8twIq2dhSJmuorYVVFwb11FpojwBUPH2+7Q
+IbMnYNyotjQ8oFjknrZ1ikLpYOwz/020gJY/ZRUw8TSshkyPmhkpj8IqMxhdEtI
ZqNWaxIMygpEKybkxJmvemLxMtiFjWAQ/v8jX8ZKq86u607dxjVTNzh65DlwbEiH
DSz3r1FlSc1dxAjCRW5gXhceA50ASji1QvCfF70XGrbQXpA8Q/UpINdFY3lr48Pa
ruMrNZXbJXLmwOyNrWMVZ8HQZXcVXfR8/HOQ/XN7fiiOE2+/UcnZuKzt+hq4aDJN
PBeqVka/aYF4g5aOCeLO+MoJxGlJZyUaI2gx8Z7ht3D2cmy63ffKoxwAQ8BNjfaC
fg8nKeMUEJVtNhOvCCNgGCYuKc1jB8tlosn5ESXzGkDOeYnyKwGlhAWku1flu8WX
q0bfy6t/sqUV7f09LjYUwl3YW62q0od7c0tSZJ/l6ECi7VWqVJ3UFSSUyhjtObMa
i9mDRCIIdWzqGdjWRWhm0gVmIkKNwXc7sP/aOzGAvxFcB5W1BnDqafp9KOB3d1/b
zLHXgaklNAg+MCs7fPQTnT+TVhqyHnXymr3Asf9Jz8vJ2d0EIwacmQUpaH1JlLbI
7hblrWrhNTlJE3i7loNI6zQj9uFEiIsaXNk9xyFtdFf7Wqeccw5skoSYgarOE6vV
OqosfH7jYrChPg97IIoXJM65i8Yry4FwZUXS3BQ9w07AbZXnMn3gdKBP/CsG9jk3
Hvs2+LWQnWAjGMoKj0VOUGs70E++jRWuburkmma4Pbe1HZk+gAhBVc1m1ubhKLdU
dmBYZvcSb3OxRZZiw50pRyv9nZ2dCJfGHrhm+ALamwLBwEqQzDl6Yds2yVFKNsbV
m8+rTUbv/Uk+CwC9HvLzyTjv8psX5TYg8faYY46bAk70vNu/8C3KivyCiCNe74fb
5O2pbYnwEqsAVwiVajUcDpNNH7vNsb32tO6Pqz9FsW8Nr/B/IaKRQZn1ZbGwvn47
awEpqeDoJJMn+NpxV8x+wTY3+lYiZopm2LgBM67Wzq8iNmZXfFpWKwR0WBVvmOiL
MvoEelE9tVBlEREMPe7H/cNFmXf5ff6bB6fzTXaaOfVzG8NevasUbhB/RVMQksnW
rOEgP0fhvQEuui6LxU0/P+nEz6ol0lEC5A+TgJ/JROdpsX0wgl4kTrfUhOk2zR+I
Hl5Yho5nbJsKS2IljHUPPHZd5390GRjIEduuIvC2FEBJ000BDCFOxxVguJtl2fr4
NYTTHeM5KA1oq79hgD/Z7yPwbMSwm1CPgyykFhIwu90wsWKEJgwaRXImgpHdhk3O
PJL1q++MxHi5kHmktHaTI+UQlF2Ju1aJY0e4Y2kWBtbXO85xuox0Jds9F4wJpBm0
mdPk4MztbWFfzJNdqvH5xRPlDAAxjSx5lzuZFB5y9hjz8mWUrBVTaVy6iWJ0SYvz
q4Iow+F9VmofYL+lWld2vVYF99osVTvPpT6aVs013c7O1R9eiEmlINQySD9UTs8j
WarU7rfaGCuDltN9e5RjivkDfrKdQfGyhr3VJei/ox50ywYPeYSfufWtUiOCSpiA
UCQbwBVRGG+To+iIpWSUOSt824fswZFtgSARy0fMrzkR/9OGkanu/uhysp+Se4Rw
44o7TrJ46gExUs1BUX2cdrQUhraJKPjfzZQL/KaaqI6WrUpweLDC1Q/pc70EIT9r
44OzHsIyGQBzLc1jn8ED9j7eRBomhY5TwILQsWg43xzUnIVoqx09F9gJry+9IgFi
qxkkf6iDmAC2fcKqH6C6pyvPR4gob+L3Lqcak6WxtLPJn9wdB/hfoy8++iVwQkTL
l/9UkAIr/4QvZSFmGhRaVZLnQ5yqDU2cOrigoSRfX+VZe3dtF4eSvg+3Tokxdnh3
XZrxDhoqXwxV+z9r6DohoqR7StTVJ9VKFb782+AjcYVHhm+rCp5fTNdQr9KkdpsT
TA+RrPRoAn+iwbwNdjnxbicZqfgBgflZ6AdzQT7SoUHmeBeWQuheyIZ57o+9z/dd
wswimcQ5/WeYr+uLTQWI6LXsPJA2H2vtfrWCqvHqpngEZKW7Ms38i0J05zXoZUhN
6p+02o8CwaWP7P/8EWc6BL1dlOxebQ+WtglEAjTt48Aad75wRhCVpGmk6miSFQYr
rPbjgE4lJrzTVr9b4nZ6yfyaXOMgno/p2bm4i7p1CniS3arbltp7IICGvJEjIlA4
cS3Nu57ZeZO+qqv7gYS8vozE/HP8EtlrxQv2E+qJIYX8k1Q49eckk0Jv2xQGwGKs
mk/rP61cyp7pdoBYpZ8gYxwqb2O+xzo6IwtKO+nm/0VMrKJuSpzpdZrx9vKZjRNd
Yg4pWxhln80/tQqE9zf8HUKOBFsu8wCmVCyUeXSFdh56ovns1EV95jymCunPUw0L
t74TpNmWqis3B18goZKglci5Sv5wMuEM7b49rL+FOUxvT4AKnPRqDSBwEkWekBb5
bW4hE+eJIVe+n/oK0tyLzab/8dMLYGIfKvlZDgMocF8i/rYXVTvtaX3Jhu13X9CV
iT8BGcs6Bc3NOqSyNhmHT8h0unkubJPtOWPIQYLeoxUMIcYubgKRq1Q4SMeOVrPN
xN+K7coTTDweUqCTaxXtdxW7gYhduMIiJMbYkNWNZSoPGZPrVGfIH8mJdMqPuDrb
wfeQ79ZpFYh4AcSM+U8SZFEmDyglay5PfcsHuQFRDI4q5/SFUv7YV0gGz5poTGlC
pOMmrJJbqCCjLZJCkxlXjyap2r4bIcDA38HLgK8Jlc58h4wwiheqGyVeRndgPtkz
ADSuSHU2AhKIxmEkuGL0xQic3z5yrzDXLej19iBcABVmaGf3ksU+XExQAyUzbfcH
nA6GneSoBrcqBiCWLg93MDWjJq9bqYH2hSJoMYGX9mi6Qzd8zpFPveRNVwXrvM7Z
1nllESoFWrxADECUxmZXkAwSmBtNGjOEY3ndT4J/dIGVSM0uRRwODBLfuH6Bx8M9
iOM1gO1+V35aPFycE9T02v13CONdncNc+Z9IGBgQ9FkMYmJL50d0EVOqNnLTOQb3
Fq4QCgM1gMvqF4dCi/WqyQ///vAhuK+76wz9GfV9pkdNIAJO5+V1giccievSPtFJ
zkfTjLheLuOHEFhNgZRbLatFD6CVvNGnNfaPEIvfifDIqzddQo9rsVThGkXSMJDM
XgtXt+gXNehQHaQp9tOGLEyQBBkl8Mc+EHzi9RWeqINPhhsB16JNKD4dfmq+gKcb
IxRuGrzoT8Am7kZsHGvXZlf1w/z/F15/ngyPswr8Dvm1Cv0aHj1Kr6cwIa5PG1i1
1JmUormzh83Pt9KkoeYgENcYApK4TnUiws9mcTfyTBa9+uAg5DoH3I4S29wXF1TS
7zBce82PmhfpO/51N8yAEluX3RkB3eZTCqRAB46ldGQd6wg83i0WJmJUs6XjMDJU
sPoudjGAskzJ1VDAOxOyoDoNbZJbDIctcLK6NTfyH+1KH2kkRZ6LsdIh1LjrlSE8
UWRJexEoHJB1gLhBdkiF2yuk8NLaJAU98pvhqVBNo3US2mJ2fPfcuna1f3tA5tfN
HLnZtl/zdftD4YnQWohMizgcDaEHknW/B8hfDGN/GJ52bvOnQo7Mj+p40ddANSGR
pd5DqNXaQ3ApdQYwbbLKfJ+s4DT31p3oB2GIIIHz+Q5K8wug878nEUYvc6SchPN2
7VzHdeQfRjp8dYcGqd5zCOOSxPVKpcWKPzYzldJeY8wb5Ag8utJO0Rq5N8bFgmff
21su4ZmHON/vmYHNsJc70WXwvqwJ/BhAqCEgIjcbRiAtTxKhm6eVFtNi/YVyV0Dr
o/Zs61pkXLuGtIJaKrEGd6syxHQexa/ROZvRnYxftr+MaPfv+QuOP01LYxU5cZu0
Y0LKqU/EoKwVw1ukHumeXakStFJ8gs48LjeJHdJsl7NljknTLvpn29ndN9kfmdvW
CIFi3JSQ4kwzHqURInSzxuP+MPDw/rLgLm9BbTq1wO3jVzYciYfPV6ufqtrNcgMW
S7cCh6/Sfxmupfr0AE5m9LNYnpTmbQwrI2L2hCTlDkCUBr8tY4SOo4F1BuubT2vS
pf3JvOobEGh+XujVND0uxn6T9kE7BOiAy2renEcGLpFO4nzeVfP836t8os53PBxB
rwkGgbrROKqhhDWRN5rhIJQS5G2XbWjvZySWOCZKdn2wadqgrKGGJqTN/1z1oBTy
sRrmX5cJoDBHgUWbySEVQDqXZ3LcmqovZCWKVrAi0KgQfh32+WtPn9gQqXSge4qd
L9u28u68kjTxZio7K1Y2dISJFxSOeDa5HT4jjwSdTUVvw1bqMrmrRaTVQsEj4jbC
0NUpFV2CDy7tSvKbaN2LbQ6uYuYR+DPgmov6gyyYAuOhRIYFOlP1gbExI51AZOu+
Xh2Bqc50ATyEeRPsL5jAByPhMVC2DlPcheAu4zrvpigMrfpc8XuUngWF7qrIwWig
gB6FWK21KDvhMnD0kOSmE7e2JkmmfGP1Xf+LthzwlqS9qcDhKqTpgCLDSeo6L7ER
prEKFR4wXq7PMCXTl+m/XsoE5P1bsq+bF7srSqj4JWqmGTS4OZuBvt89GmLos+z2
y2JkQytYgmWxg0m3WSRTIiNdYnATNrqo3mYw3zu1Nr/8Cb3chHi7NDNYVaHW6YE9
SSQ9B7cy6N9MMAYE3uwGshGlrejy+175GooSQzyQY8kDpMgf4vL93XARKoZ3L0bL
nKceGITNpdlya64Dt9jalhLLKPIvGAzxUKSjELdqsnDLn1LzWKWV2qgcQtn+z93N
qZY0SZlmsyYtp/+g2dEhaoeH0/m9BsroFxz04pLewmYB6PbIAwVa3f9NAs33NZfM
jXXGAYVBXU40qsSyN3BTxHNh7Oo2BWZ3Xx7pM7nUzTkMiV6YnNonk4H4YhnzPkxL
QUyNaAwpIoDLULQ4hjP/mcIOTYX648eZTOIAITQ/Fp4T4tLUcJs+JVnLsneacGl5
FZhjy2X8MPT2r3BY+llTUe5FaBT5rlTl+gnRuJiSuCVIwhl8IzdWeHgtoIzB04Eg
xbPJs6aY+a5lOme2fSvmFIMgOuTI+t5In2ZWmo/QczHZcDU+RXhT2XU4ykb+lL/i
QCrmtxJEEZ8+MSbsDKGiqf4CnKLgIR7QwNshl5aP2KpvaHVK8DrZgYHpemQbEWry
W8Y6dADQfDZ2aHlC+pe+o4VAT01w5Rza/ythrcbQvLU2GQV26GTTlwZe0cpQj3MO
vICNg0j5Xb9wYKRwhl1KFNDlE3+daEgTDDJ+JpqwInOdpddRoUggg4lcpcYtavzD
r8YNKRDCyPGnsR4xmq+e4M1RsT/NKVPkau6Cv1WEVS3/o/kJBsyo7REhq7SdRFxC
TZKma797IsNooMOz23LPXnoYrRGlPJm6M7cxQWGtA5Y8CM2DVEQVr9d7w1MFELDI
Z0X9HDlwZtfkoqq+/dqafMwy/18ESoic9jySeNwdL0+jk60EC4UAdVSoFiB3tvVS
OaSIg2wzPXH2+BxFAi8xmO4nLzWucsrwY/RxW2jaOqJ8IdLrx381bV3vhdoNg0oo
xg17dB+Pp4rurVyRBVSyvQ/Z9dor9E/t/UW0lB/C0u9LUhp+03AFLdKG0BryppF+
IOCSt44V8aZmQ+upVzb0r3EzZPAUvyu9e3xkWcsxw3eHIC0yPLxQOgeKkc7NAbzX
NDZjH/DM4CpJ9XTnbX6uzrNSBKfU4LqS1KjMLkQu3sZ5U9SlYTWhhbzJGvUonpEw
QxVuwXdCQmOd/F0NElBalwTD8lqRDnDmyxWg6w9g6xvnd35OivqtK2Plqn/KP6yN
vT7CaGTTxJh2hRF6mhDp7chjcyqIHhMWcYsAECRQRJaOsDnnwQLCiU3Hh9UQpAze
OT98Oo/8AvAxtYkOzDMhWiK5ZkwjA1tNq0OMFiMSGyrYAtyVXM5KpNy8Jd7OX67G
OE7CDjX0goR8qM0FyfSzU5Rj9WrsNujxw00KlStbJI68yxXF68bINDDo2yc+e1nR
omC1MO/7xaF81Trb+4CFmJeKYeM1wPYARPs3sJQlFVCOcNaPummnrTm8AyJBrArq
7ccBC/kv4/9DTyaKEW9rcHrZqEVkZunzxCj8BwxH/RthDOIQfhGBvTEx3T8/v1+3
SmW28YeZKp1DSDl8bJ+8y+la4Boo24REDo4izCoPIVAJFWFSz97vM9z9+g/VAZMH
FX8fVlhjqi5P8UTRVAVqyBAHDzhIyrPVWcDw64NW6vgq7RET+6TDwbsSsbzGUIN+
PXsHTA0+GExqUrE3cnA51yH70fb7xnNW8A7FgmlJnHcn/IGn3FkiDkBYR+il78+o
3nmS6MeblyuWg9iO442geqTrl3ixumiOcdzlr45WLrbo/sbDpDdGpOd/iz8a0JHb
GI8tDeJ86YOZevI4rqpdhMien9bB6d5JNWvtQ2pYGrdphKwAe/msy2rfx3sqWuE2
Q1aeTweJO3PwcyiBWQ0QcFAao6d0Er0JpDdPZ15ShyL8kWtWIs+n4y0sQ1yNgjCM
+PAHe5KF/o/Su0nZl/+EPC1vHdZ6de0ZKXEtxn2BIJ1266OVJlRwzF0AWPxUS/7r
Fz8bfkfj7M6tMWWHb76Sxj8KZCL64Ov6Oburc7/5iE6Gile1edeuVvpSBSIiBTvB
nj0zrx3sFGPvzhEexdMKE2o8TvEe+iJ1JIpeugJ3XQU9Sk8SKip2ruk2PtL55UZ/
+VevrivYB2dhcQCG2oM6M9TZmxWeN497VJdiDzONN4q6sX3lSdGrskwKQCISVi/d
ZXc9J5LSVVEKSjxCdvfdoxuc3JCO9P41rKiOwsx2nyQ18ebY3aoJszB9j6Nypbqy
UTLukdidqrBPs4/B0h2WR4GnBDT9Lx+kpukap/YjRlTgOdq78cLb6bpiSMVNDEdd
+iWN01gN3VGEoi2bYezCUvkgJs/rBBCxUNTA6+Q2zb3lZbBhYRzKBrOD31LEvEKN
2QU57mT2dGrG+qnSK7LO3NFlQMuoTDi+Ut56IFKpTIGT5Zr9URyxgvL5rvFegIXq
qUndv2vrNpaNxw7HeCiveNSpmXRbYz+a2NdiGm0mzMNjqSBd7GlLBM39lt4K0uX2
MlWROfNJjXbWgvN2NiNX8JiKeF9tvOGia1KM01LRXvUfptmGvqJDJsp9ghpLOG5C
0lhbDJGfcjstV7q/HRqDSMNEmjTjmoqhYt+l0lzCWXEri3fT4hhT1+c267Tyhf4q
Uv4Bmi5caFwzWjVKshjRNbDJPnZD6Vu/IGaP//xICwqxh2Kb6tdHe3MHJwneZPYi
TibYE5gsnVAHyKtSGDmbQgmcBItoLrtwyFU0RMtc6cj4Z7TRRLp3tIphDYP4Si+V
QYhgQAgrgt5esWStpGCS/qsMOrZa0eGwCquEs66dQEZc+hilAIzpCxWVXdTOPlR1
Sd5qg2QPYUT1D0BEhDLNoRTQyv+QB9r3utZq3T0bGTtnBVZ9p+jBk4TIol0IKujK
yRApz7FskpUaPdp2F96GoX8HY4OyEq7fcdOH5toq8//GQSCd2UlIFzIDBfRq8tbF
ochm3xCa6jfQMFlPTNRv68GZx+fu60jKBBcvthA7f0RKPKG05XGdAFgNBkLAlQUD
X34Vf5Q9qq5UqxCFYEZc6J8/35j+DFdcFZTqZ+d99lpsQauUfBjtI/NeY2KiVrep
Odqa+HZ7nIctLCIApPcCNiVYxD5Ic8QlJbR540J8wBRe54kqUx1VKrajMAYRVtfu
ifCzh+lF8ds/3vItRjJ0hZl4JYJ5pZ1VsQKVFfhY/eRX7xdWNG188tynTEeOhRLN
5ZazawraQx3LM6NaRegpQqymULCtj415A4lAOlVmA9G4rJBIYQHryH18glpE74V4
bvikV+kLLThKx7X0s9VryxYrzW3RjYeMfOjrY5gP6wlOcRKJzi9Sm6Vk/BqOs9rO
lzrHmrlCw1uF+Wp0AP03soqkZNwhKIl7UfnVtvxJtzOeQr9l51v9bFA7K+wcR6d4
r71db/SuhYaAAHkV54ZQ56Vm9uovfJeGYDsp42J2SDiYdVyjTbLf3RzE3OoPiZPj
CrecZFX42bBn7S3wqsY3koVI2tXwcAd7u3a5dnKhlfw/IKpwk3tB4YXByGt2CEW+
Wjot22ho6Ru/zesYUhTkxNwq7vybeMhAWDziZckDsaRv3C36aGCJW1YQw+mV+4BT
lTnS/fDnWr641WCecTlyzYZjFMEaWaEGOg4Dq2f0nFcDlNr3W65NeHgTClKD3BGx
MxmFdi9Q5cF5xK/l8vxWchx6+lyTqixDmx+ZriFabHaHFYq3q+2Yl8TiTuLvUJbi
U9zknVmyjO5EAHWSU6eCpXUUG8PUXTis+KwuGMKK7g8Gsjppr94ODqAnLEsmS9po
0BnP2cVIC6AdH+aA4XVGCWtely+F3wdwq3E8XJIscrrbuWVWmUIGE794WsXjqk69
UgYhJ7Ds9wbhuSMEdUUcBte0XJNRfAU7ea2GwzTHWiywz4uHVUqc0prxB9GCNrUo
twki2Q1wrkWzjI0MjCEKVUdw6MgghW1JKtYrHDHWVwq0p6F+r0f/xwgsF13yW8WF
xgMCAbW8n0todFGxebzx+rNIyD5zDtWQJqZT8zERp68OvyHPHQqfCTNDZOD8/YbE
uMUAv9v3iFrCrPwkwBpyTa/HHPeFt/cYlQAuLmfmVqqt+dlytaX+us3W+y0JTh+z
IblvhkY8tTnNNJW/P5CugxS5ExAOcAo4exzhc2S15hKSOsXavCeNz7a829f2ITX4
M5dbyPWcOmROFoEJcXgFAWOQl8C6rj5w3XR3WdpXcvfChY2z2iPYvY1dFGDFls4j
Oh+/4h9C2FmAxYiM6LjSuqhGZFRQC2QLvakVGvR0HPP8RyJXAktL/8cbl5UTgwqJ
sXhqh/5mtEFyHhiMbv/o9mI/3a9NPAQR3j146kYvfwvcZ5mASxAGTi6SLD9BbQzQ
MYlts9rsLwEPvQEWdS+ir8sZeCNo6GO8+xHGNno5ESy/35yw8epgZpHd7FB1bKF1
RiRVJAgUnVTELbel8Qj7j5iB8jmgf9aIL5BL37oxrsV62hy62fxzcXrOrP0upC2x
yXuoTrDBcxScZ5x0l6SaGegZlEWCSf15ftmIoBkck9i3rx0EbcuGMfmkbwyOHV22
btGkRga057Z6z5o1yXq/4cahGOt/PSWUebWWXVKxfk9GJtiGLJztU7ndvibvtRxa
lh0AuAL5jkHL+z0bi7xAT8VtvxRj2TeTI78duV7/GWNoY8Fzjx2g0d0ulW/QMpdB
w4UtncLQSxK7kZbpF9qu3/u02QUNDoOaurDnTh/BkSEQ8Y5/U5xRlODufXEAS1lJ
87+2UhqV0M6LCs1s7X6J8uyHE0B+/D3xttedUJXQ4DsmlMCIbatGRFdWNy+Qq2uI
fITN1Cdji0t7q72mONvth7F63b/kHbHj2d6oWpgaRrWdHJykdyAultZ6I7qCZGtN
UrelwFcbohrEaDVgooADkIzkOigUnnddxeBWH/YwIDko0Vj5pXHutHgoXp9R8/jy
18Fm7G+MSJwLR6DsRDVUbiQyzJIB0/Toy5pJGRexwiUdi1zGfLZJEBPKp9L88SXt
XO3iI38QspC+/hk8g1d0KX/xtGbpKD1Rl9U46gXAJ1WAOARvxrBGdKujamINTi4h
sA7929aBjwLZgeyz7uoUEFo65ZmFbDjNerQmpszYFQXZfHNLB8wEYVJWIgUxIIRU
yrBsiig/E1Wt02Y1tPAc01sIJkFIQEzeDdX9Bz5gXfMTKzF7LCTCQU1lKNZCnt6w
d8yAZNXw9Teza8YLdgE1mIWZkSL+3rZd9GkPXpdT+dZhLioeeXWprXZ8XkXryfJX
NvtPiyGRL3LQLF7SL82/0r4LFrDBohncgVuUHn9BueioWVchXAbyb98DgBgieHwx
vjpWvcZ9Qot90lhLKqHHT5qlvlsrObwROtQNZ3ms4rrOCHfMyzUT53kXuVx1fMcv
JfpCP5FNbMf7afGGvF9XQnSNSNcvUIRabYKFzCGg92u3ckb1dHaYVjX+UBYe/MhY
sBoyzNqbq8K9jfTN8pQJ/sXRk2Bay1O5o+Z7snJ55BeD/GM/6pSRp/thAHoD3kN8
6PRPUIH8ScosqULeFlgXtkHjGec6pdqRu5UhcAt6WdPvWUiWV4WKX6wgAjCvDJIV
//jst532ncwbXNz1koU2HohMp85qQ+MEW8xHz/wGdJNHhCX5F4UDuUFiIcCskxzC
E0mZohkpSbsirdLX4ychT2qqU/7+C43DpGZqw28EFd6n97bIjIHksE5LjpqMIXSZ
NR6zJ31okIPkUOMEnEGgWnn8c9tBM1uRnoBnFrB+athFRytC7v54XsRXqYSMKVXp
zCjLIfagcB9/mrOlrYHNQWazr0WobtKXrsgsZ5gH1stTetDgfbLR2zg4iu/NFI+Y
XHGhGDO9Xsg1HiseePfnhHS7CU3gLgvDmBJsTgRLzOa5RVM1xds8O4fACj1jSWBD
M+TRSIYpvtReOnF6mDaMyGUSqIU0rTPstziN+IQ1eHddKe+qraZaLl31UtpwOur+
vfqwvMWsI5S8y81p5XlN5+k4qEk52bnauayZFaX4z3iqU72hJdJqQD9Lhtx3qteW
T/8H31UyglixcOxhDqhzdbiMqmrmt1NFawOTepe4ysJpIIi99eel/zthxLAoXLyk
BZ02vt/ObEqMiHYGGijGZNqfi6nW8K5SrZNyM/NAPS/VZcRgLkSNQl9YR7jEuoz0
lz6+GuiNIqUG9FV3AiJVEhyM6f8mDq7Gw+ws2FaJMHXljDtHE44DgJixNZKfojFF
fVyAssqyrpU3lSXCieR4N6c2+QWo47e6fXpG9cLdbu86r7vwxt/oGUuVFmdepTi9
amr/L5KKT6J4t2t1fqfR8uDldoYb4wfWnBkEVpjBaaGibQ4y861SsYXQFJ7YM6yp
EM+WfZF0kF/6WcPKzszj4dBl6S9nlEjFpaCsaA7mstmg2XbxgbZKpj+bQ/LkDaI/
bvk4Q3HHmIJRb6nFqYBoT1jc05ZZLQ4IcbE54v1yN0o9v18Tbso5D4OO7bNOQqjP
m60S4KJUiUJ0dpl/kNyNbe6x+tQWbfrmXliGcXxYiFY+pv7MFCta7FBgrKGXBhM7
KngWOR2s+BfivNcmCwmmUmFhdTmvez7mBoA9PeBKXT8ec/twQPUf6VJnUZ5B+a3m
OqEZFgaDlhzdhP0PsQXC7WuA3PZpPBXCariwHrOqbjEH2JL9AAWzlP97YgVwVfWj
32IpT9SEnu6I8VYvUCY3BNDplTmPi9IP2vH1O6wpU2zKwNCxkQwfNdPR+uAfHu5W
em+p05egofws5/F9avipuRiZ5b8MMwoC0/aUKmGpuFKP0Qgq2xrDlwEeauY1ev60
wE33fg9SK+1QPx7/vhrWySocnjBuG7ElGzk1Nv1BxOLeMX/BLBJyn6QxK8khr/L6
nlK3iVhLsw8g/Yba0W0+AwbOks2QFrdw/IuC3N0xOvsSXR8IgBDYfhoAL3af+PLg
VpseelMDPSdMK6Yst/v4EagzTrBmv6zfjt82L5Ct/WPGU2s3VR/LcNSa2m0+qLyT
Z9fBapul+Ry3Fivq8tPFXkV6kuWAPV6f5uroTHG0xP4w4A1p5H3UhCBbceeEoEIy
86vQiWyt/bvl1r163rvrwXi+YiT+S/MzRPqV6qMu+vXqOgXx6Fo8bhJZwbU4ZppP
yU70T00jJ+P4ZpdcGErtol1XqZllthx+oSztDy4cSmK9uDrKnulhosHSRqIapDJ1
vDiMXKggBL7pZhhFiVHiT6gG5uuQr9YpvtcG/8Uzq2q+Li92Nc2VMTTdQwLxPRYx
Vw2mzTgdJuBq0sm/vIgdM9JkEhFnFd4McYtoqd/k89LrlRY/kq/6nsPN+rejBUez
n4FmTuByRYZW13vY+su9GkTp/fGLTOyxT7M6LCrLYZtsS4n11eHQ8ZG4sj8u7R2z
CuphoALnbVzkLq/ajfuoDjHsmjOTjqTpjlNwh8F4nKbZ1BYQxt+qL/Fhijj5X7gT
QC5jw3oD6CCoyhf7urYBvR2hoiJRuta43IKc2J3nRzYx34EXzf0vTvEEdqaYIw8Y
aUTWOzFAGf5FO+CvEDdpDFPpmVbJNtBEIlcq+l9730ZEB6FTPLdgT1uQDJW069Hn
rwT7qPjI5lnDKdgmLqgaTXUC89WwvNIhgIre7LIINSv87Mpnnye7jLagFeIXh5+O
WHv/TJlqk9vrBv7MWIXifjUUSe/18tKfj5+IpWnAO780Kt4UXChPLwvhQ+4qqKny
Ttjz5qIz6JVirTBUe/f2AwFyYa+loZJJ53Fbn1N77O7aTbhdQYbLszhVSihL/hKM
B+aHCza8tG4962imBCYclanuPgMu+U+fkuuDZuQDcKwISB3fYzvxZSPMUcPoFhRQ
9O+KVJRgwx8nA/FR9p+Ps6HIAjAuSRewCF5dOVz22fP929ylr3Epb00IGh5jbtU6
YDUhZwCc3DFSCruAMj2xePEO0O9kyJpMA7DRkRdGiXILq5w2K2mf0OwrXQrFD8v6
WxFu2HQ+PXUX35rpwzJ755iNVF5e3GRCp/0Y5yiugrk16qsrjovI8JlUzshUOBww
ZIm5XdLxhc9wcijDCOACkc/tRreus+Nd5x/MlPuBy6dVZQ/GlBL/Hsu+fW2XyxoZ
IW1p2Wm9WvnXOgdEKq5zlOO7/YapBW5rd+TsBNd5yTghLN2YNp0nU3KysWQdrMYG
Dh0A14ShRRQa+dUlLB6WhJIbc8TIcR/EXSsLgqVh+8FRkyD3NTeBdwNtNJh90O+q
PZMpDHepjy58JMfGtdFHrAYv5Hq5Dol0RxIpVrcWbsIyU2sw32i2e3jo4ebxvo7w
IT4oW1YDpOF2R/718oAPvumFDwxau9I8kHATMsiWez3qZzDNxrug05Ia1ikZvZxB
Pz/kNRMOqF0zf6awfqJRWI/vOUMdAs8U35jh1TdoY/ofPMVPrlYyQRX2MfEVDRh7
8euWLFlUZZkUVsiA+ZjL5+XGADI/IGqHYa+TIwiYeZEE3q4kvCR/rx+MkWLaZKXG
JB1KMuZEX4IuKUBfMm3lhTRD+gcfuRCiD8gRfX/4ZpyxwP9rwnvBKfX2G+N66LOV
a/kDTKsP3lyoc4lURZLWbMxAyG2tIdDO0urV9rbO0ykiuwU68FcJGkHXzOhGLKNN
v6JvPBo6VtwJ0lY36LfYHJ6ZD7CfxsX3Zj/k//R/2EpGJKuudUU9QDXHmptzbh7k
k/VfmLwU8W0S+qowhpluGK/LXrmIBWJWYD+rWLbyVBliflHbRd22nn5oU9NLjpEf
lK2fZNUgemDUEYpvY3A/WCCva1Ym719bMXNSDai5dUsgarIhWC0b9vi3sulHKMcA
+dT0H3Hx+LdR83MVhX314/fNI3KQQh2KZ7/l7simtwIeYWjiKAZYeUYvvJR8Y3Wv
QLgqbNLyqna1NBH6d4+R0Q68fLbdUBdBCu/EdrTjM/cPZmltP70jod5lPmGEsJXJ
0DfbIS4z5QLI0NS/kwCrVKtv289+5+OVyKU0rsaZVMu1dpxym/k3Gi9E57+dBlRO
iQ0HDCFGlVUyE3dmAfPiE9sENRM2RM+jCbuYL8Bq1H2DgQ8NWO64AMkAJBhv2Ymp
2WEAtJg1PoarERargwnEP/vtwhZTaHconChklWynBjC2Ljf4KjfmxpaNhptmtLS6
HLxCkQl/aCGoWpA++Uv87kpKPBy6Lp3PQeihg8AcRvHW9PGxtWgtY1amqGtjZ+9U
ygerrx1GoujXwe+gGxxkmI/FnRLvVNVMRXlbUVEOiqkiIxtnTga1m6dg4+quTJUE
aOFW5qpbHWnBOH/RM4QJ0dL5WctRibp/zIGiBaO978Kr3RW3R09CGjExm6G01NdM
5LL6nEiofBTbaKlXUuUyg2fpFQtmJ3lyu5dUlWE9juS8FITaObQSH6Nnwl25uDNw
RB/Sg65DuysqVgjGCP3UA2yIvrxllYMmbHQPanvkuIO0cCxbLz3sAdyg7xEKQhvM
N2NABwCWXObEoM6p/iWY/K/J7z3GPnVv2SZeA9n5Hbk=
`pragma protect end_protected
