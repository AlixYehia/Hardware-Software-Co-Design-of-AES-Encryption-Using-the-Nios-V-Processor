// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
oa92VqD2Plhq2EnNFG27b0y0QtRqX725DvksHsJOPIMt86UfYnb4HbdBUm4xHIp9q1eeg91hQa2t
CQ3nvyDk71CVxIA131x0/ujNhII5taFSmc/A/bBMzJ2epoxo87IxY6bHh/h1W1IsG0Xr5CEF0flX
L0OXC5SHgsx+XRAnnCWGbyfovQRW9E6wL4CFOHXBwopBNaDdBd4wnvJ/4g8boFCHIMtrDzLOOpTj
5QLM/+e6qVficHoq5CoGVrbYsscx/tPLskFLiLBDjk0NwouYTNjDxMkDCxErNaRqv8XNYlob/PXe
JtjgG2bEF+RCQKvVd1PE5ayEM+vIMqY3z4uoKw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6352)
hJCtbcZ7vwheiHKqqSrxsbAAJ7eAuSWg1o56X9K0wy7/HtSSd5QURj+FgebZVFiVKpUfbAY1YqkF
Uloyiqio2g5Yw/p7EWReMjEgtQzKaqybpTQt5DrCLZTFqnAaCls0y9Pez73HSjDJ5OgyQAnog9DA
V84LtzdkrOueTP+a4hsaUzZ5QrPA9dNDJ1KDGfxWaFPjHMI2PDQ0aA0sEetbHcHC9Z/8TwuTk7RZ
l+1NtlkJVbC4CvE59n/fGOTA8/tIbN407L/t3lhDZxb85k4YOwdS6J8Bhvk0iOpSYF83nxZX3JuU
MqwlvL9cjZ2UcBtbegXplwoeHCLdCRtxju5CEEDbQ3NOHrr82ESsqwJMjEY81qjMgaSe/EnqSxQo
J6nL+b6BxNLo+m2mJC1mWtbINOrqBU+RFiMlwCx35XQrdckW91Mg+Za1XEWzV0Qpw1ebAQf5tJlq
/V6DeLhks1GJS+msU98soBaD00/T+k1raVbFUgbxNLxM6kO66BwyW4oQ7e2FeEXPFrQ6BGdWMNy6
OPgsaLVAbJ+oTCJz4dpmua8L3wanmYkBOuMZneZapDxlkQzYgkaOfThBBIrGGCUAq0ia3chG6ArM
gEURgPQqlouthMGYsUIE5T3a4bvx5nAmENgiADuTbX0BB4jU1l6QsXK7v5C+BLx9FXveh7kezfuI
BKTzucIbVNvastUvfqxB4sV/1j69P1hUdXb+6uBG08GhCPGCMWxdHl7WQvnBEfgQjBZOFParz70j
xGNLI9mTAiMFJm3v50898X7ppRtwADIPrYdEnJ/m/Wk64iSIrgR0oFi/F4WMc5++cMnp8pNwt0+j
9F86m748Xl0ZpaG42Jgp+p5zbAT9yeYhzHn1YRBwvtQXToMrDYEyw3wpQgtoSx6SIPouNz8j1WHw
ieTf+gGugnbz75h7gfTICvMF20WSYeXEKCzRObaqMFd77AlNx4LfnMtloIGTfvmD5k3fBpRqfPFD
u8/eW3o30SLHmbT7q4hsFR5cfS3FljIYHPZrHKNCOntTjGxzDFE9jAfXdaQm/hyfS5LtoIGp2qhr
0PALe9cAi+g6ZXuIHiCWi0e4QlO3uleCOClJbwvKVqNaoaq9WaxCBvpNGrprxe9HS6wUiR7CbJ2Z
O+H8Xd4JrwGTIJU1ajNEzOSr1NL8YHcuYUqPP5Uea7XVkmR90SduDGlnBKjWGFterz0D9xNE+hM9
XbAHP1TYdd4JPGXp1ZmPLUPgwsQJ+X4Vd2DBPpq16ofoXuvEXElnHpTTWH4UsBPJjQYRLt+KLXMg
TfYfrTCDxgJRJXsXd5zgMbr5RwEdmnkwiPyI53ZhKaiSHlWrC07TobGOm/vdyym3wdwist1qvAgl
KU0fGfZyL7yk8mCBXH2PXeixWDzjZb+ndD9tUXG5qq92ndPKP7o5LT7tJQXcYLaM5MKzUSWUvZgR
QoafsOIb3U1HGW3JTj0G6vrwkyQfi0Bkpnnid5N0lVY7XJRJgj34dA53Cjtlr/gtHYyp/sTpk7h+
7FtoPp/hTZo1vPvdes6AR/gejBsQ45sXcfS33NiF00zZX+0TcGCtK8KQDpvfGq+03Mlr9DqUPa0e
0yXTU9X3EjMgIIwCjf8ofJYpRCz0an3hubEv1CCzLP5yeZ8fKa2YSxkCdaf0A19KfoZqQ4e2W2Px
X++0ie1WSC6nHQG8bZjPsErKEFFjAaWS3pz5WHetibO8cmLLI+zNQMHob6wE75dpLMNl90V64lgk
I6IS4/6Qwss7smHRaqBe8WxegyStf2Uo9FdUI4JLpBBR7HEiCLSG29Edl+v+yhtto4w7rcm6R57a
JB+ymZ67p8GkAjqsONpuV8ql9Y9fnZrTeAEM1mCkQ1IKuMBZhciamOU2LSPgD1XBF+VMeGp2OGCu
Q6FWVS/p0Ekzuq5rvsA25paua2oKzjL2eED6Mf8u2ME8PyuP17ZbI7lISnXodEMW0B5F57CcQgrI
jXMI1a3LYrurOgqDz1KvUdA+KEXGH9Pd7zgfAce9sJqiSevr7WAtQNCENWhgF1GE6ArHDZUN4IxD
dDhgTQvi02fO44zZIOTNGn5i25GDsiquegOftgbZ6mcRBiA5d7jtBtBqsWQ1g+v4i5sgkig9cUYZ
kyjflL2C5y7eniKfLD997CsRlQgDKmnkpLn1viBiA3M3Uxm8bg2D3OPiQO1H/BKe66KHJZ+QdAqg
0Y4VGiKTMqfOBomLXFpeqSkrE+yf9c2DpZP+cGdddmZ9eRvVOoMtenL/GIJF8P8+Fiw3b8Rmh78J
eTkzo9xhuKurXtyPjQQ8DrhVlIL8SqxyCT25Nr7CjTN9Q7EgXcrBzHBxzqzX7U6iObY6bhq5BI5w
gf42xQRXJc2jHIBPIlkZwzSvGMgKJdEs4NI9aUdIAbjT5OTbefATjTB2gkfScKNsxDOBqR4dINEn
mBwpOnELN0uteNbZ8dl4jroKtBgx/iFJRgI+H7MuEnWibfsWD1ArGUB8ZAd2fCsbrGDcAwGh2HSz
6etViQrqzNhFh2UoQj7O6Udb4GxlQEPqgMGfFkwemyU1qkiM128EF/viuDD4xrlEpU3F4Sa1ngu8
44SKqnTV3VRM6xx3S1022CoAHYCVDg9wDb7C7DmXUrOqrfdcojhtWGCXV4/HKj4qvW6X58VZP+VG
9cswusBqBQU9rl0HrYzeospcXtFNSvgrw/PhdPHSL6o4nPvgW860EzB8g9oXwKMFfQPFBOvDgsot
7aqWjTvTMlro0+dIa/O95j3aE8793UeMuRMgqOKQcQydEnHTAognypOUk2EOCDC5323rcXjtNhlx
kYjBAM47jnudIFzvzK3NfelRX7q47zNjEKgPcopvUB22BFM5gMbgjMdx+95TuYxJn8hGSO8F6sR+
yYE4R5XlDWX4JIA8KrfT4zrh8xBArKbMaxfDGuwjk+p62dEcjHgLfKuVKaCbh9egGaZNq9UjO/1R
rvhjQBal4qqHL9KJYfJnTBd7MvMqeeXdDs1diCX5HJQhlQsQEsm7PFuSIjDXQRTIcXOYUlmopowz
P93UxeAIonDvQ4YerQ9jYwC1CgQXGABH6KGVcQ3zCmrf2XjkwsDhKnNzbryWVF4uxn39mheosBE/
+xUBc0ZVcCNs6RoTxFTge0yrK5OmYKQmcDdTsdykC6ZeTdcRUrf8wK/hSikuHqZ/UkLpmmNeCot5
yIBT9aPDiumDBJLTMDWQu9MYKVDrwyWr0JDOE4RsUTTduz0O+SPnnkNwVbV0ieahkf4sm+pQTUva
nyOhmbOP2eaCADIz7Bgoyg+9ZSLoqsfoWRmX5baqYrXLBMlAcrttPC8vxkDP5Gu4o3n6ZrxsLKen
9NeLD4fgAlEkcaCXwRYu+opqq+gBKtv7jQMgQDi9PJKcJwZ6l4e+Nm582vdXFQ4FSWqEjCzp/FNn
FQ4DodfIKoDvRV887xVMonqCIacQ5VNzHzJrucTjeb1e09dmCPqWX8M5r9Xa8sixJbW3jcbF8Er6
1jnFTwRrXG4rIXWuxC3DFNSv6NDT9BBvwiYjPmk5JERplFI/jAN8myMlyYmS68hS3Knwjwcb6JU8
JQJjX+khOi13L4p/8biI8pbhhqmodBZEqWMQRDPd9Aw2AjrI09FS55wLhC1zLWUStqIZirpgcNFX
rP0k4vKIqId6ljxhoQMPGHIFhvfLhUFsCWVVGWF31Ldp6KBrKMOupJysr7M8pUuS1ryepUMkVmR/
v1twLQ+NEn7ZrpWwcIHRh8SXaQP643DDORaqr3lkSW3INmuj+V8hV8iRy2IiEyoWHU4MRyQfYmzt
72QnnwNSwRHcNan+d+eek7ahLIz3jlG7j2JZCE8k0F/pERqdehEvfNBcoFPO2Z4flRtU//IUPd3Y
Gig9dKXEH8lqWTZPz/qpPbDlrgZ7cbz6ngR8E0WOWwQqLb7OF0AvVMaXwULwZu0ATrgN4+9jimXL
9uvYSna+ZCst++CKyXAtmhuiPF9dNaxODH5b11RDa8GSUZW4HYp6W9dhCBMXqsA/7meCTO4qNWs/
zuhVaOrm2jaJqAx2rb8iBpL599YRvIW8aVyAHqibYsKprHaP04FjzxKdQyPwVSSmcc7l+U851eIV
JvGth3AlV3Thl3hw5bSsH4T5WSQuhllY06ncqn8OmtEws03BCyDdYqRlpdteo23gT7+BBkPq1BD/
IglCT3SeW8z5Ol1KOInoWypKrKikNWk7YFCFy/TjsGAvueQMTBMiufc8YuxbM6/flFqv+i5P48AX
ZcDf6QkoCCgeFMVVQVZJo/CQ3667kqCTFsXSrPxmIdAqB8QhJTMYJ/kMYrmm8ccIc8ptjT8IEwLl
GpIsAJzPKuqiU1mmp0zfuG1DLz9yjl9XcJyBtJk44i4dQrmkUyhjM0n7Ac826hZF4rhMKqIByz7k
7XtBBWCyXUP5nbG56H1IFsewdQLhE8nR+92XKwzEc0rQnZs4r3uXu6LNWSY/NJsdYX2cBO6sRXgN
ACuOLcvLuuErfZadHSk+H9j4HOtFoIqqdAmzIm5DrCmliT/e2ZBUW5WxWxlcEl/zLIK1KoTUtZSG
wKfkaZkJcwBao/GuWRyTe6gEMt5KLN78n8tOtr2OTInLjkWGV8GmwTjvz9lBnlzmPkMIkiVpabe3
YKYmeVDFd790au72fi9acHokz1IyaL3pGyIkZvWJd4V7NSlYXOT6PStfvlXm3BJiQYJdYZBUBYg9
uGEHOXwFi0VIb0sRf1OjDLDZFl5KTnkvCIxyCv2RSANvTgGQELKnxaAES9CgVrzXEqNWhpbjWLVR
o9yZ0B28q/7FrlwH8WLgsZf5VvL4rzhUGqQpF+cxVJd2EegAvc2ftSvTaRqKYQ8nWc3tqydhC2zJ
m8KJdQz112enDUL6JqWDfrd7SlOWu7bcD1fRFIfAswRhiXGSNueMqBtPiawzXywxhKJJhschOl7M
ygrsA5ybwepeYmhCbuW80YCM4FZw0DmfJmnxphK6qQsuEqJ/ocTZsrZ7cTkaWprHGB90ebsohiSd
3b8KlX5lxWRvpoZYSAKgqPD3zzV7fLcxLGuWFu0ow4/4ktEO8NP7p+uwO2p8pG1Kr3MaA4K7nSd3
I1QDfd8crJl5Wt34G0H9aGg0H3NHGTsxcBLSJ1tXZrq3AEeLIY4XV1WqYRMd12DsrN44S9O4Pmdp
Siw+rZWGHrVzBBjgyaRXn+BPKUJ6vJBgHO0fHvnk8pOEChQXQyvJLFK7LlBzLkJuxOk88Q749D4z
Y+VKc1ijU8D60WMqbPqdmfBS5vVdtKpdmB1v8CL3D35NEBKeUItLhAQTsunR5oGtqHKO7ZTL8JI1
ktBDL0DbdmX6C7V1RF1lZ3zI3EUDUgNWVSNVvZKxXYtYtLhOL9/Zj3K+MB0BqDIOhl6lTsL27z6U
/WCpB4WAgLInvdLx/qkgeHld4Zz1QzHRO3TFYPPEA8FPeDSU8lgtTHPwaIM9J+ioxbNC773UpaeM
80U3+g1+IC0DiFEV076eBdSqoa7GqJqtnNz4AFRiSUM0SaLS9KL5Zzq5A0ybWtCP1ViTZhILb78j
FTY/IEEnLrZjIXmBFrvjRkBvrZUXLHwc0hkedmONA1uugx6dYgzLTLKYxrCIDJUYjTR/dLN6Tksf
InJwvdgMWbPeAl02nrjZUqOD6VANCvYOhCP9E1ZIH1TfCjdJ41lhhWVgk+tJLNSF6goJD+5CUC6h
Omg69lvLE4vbzVH1eunXX/Zr6/L2NFfXEejg2HYVaTCFQulrKOSUH54EeJNQxe1HsgSEuHgtUjlT
YGs6CZ3DGMKDu1QSJYJT3aqDr0PpAKI/Uu1ADs1nbIcWKg+hK6uaorEVw/1XzyoMsdGVz+ROaLou
Xx2/7sYVT0ONEX9SJpvILjxW5og7SN3W/0oewKIDFGqSqIed8B9Aw6HczdCa5jQKK5j4+Yj+dhio
rwESlTW5zHiEXIHaHOJd6gBVeD6zesta2g1RGN6frTj0MKuYvf4GvhJ/anCb9QMyGlxHPJ2Ilq+C
z1Oma8OM/LTnRu4a26qK3KvP/1DeXrZiEYEH95edgSWdDeNSCSFbTJLu7PrXVCy5WPHSiH4hVvT5
H23DbPit0l4x64EGZ4C7eQ/yqEyw3KHJwZEV6PXHAwRbA8z1SUcgJB2+s5Ar2qcg0Q8CNOLWhsEZ
1WZ/tX87HncI6YevBCq7/4/oMIaCet4i1YocgeQwPcvMY2DXhwukCefd+Vi2KziobWyRnPSygNYp
Yg8+nFYP409qLzPDDfKOiZdAri7NXRJ0klczM6YD9vf0BhMUnV990t6ulis1qioMgc5J3INMMRKT
xF/5e+wMf/6XkbN0hzmbMNbabj1s2JjQyTSr2InQiTC6Kq/UItFtY62Y6NWEEs2vKkfdoHPMfVOQ
zWbyHpUL+l0r7f2JF+2px3vZTuHqok0Oxlu4JfeBchzIZ0ZhxkaiPkxu2VaTq4pFMijKVJhjAsF1
zQ45IIZ7hFlf3INZRnvw43AcaisMP9GciYInlhcNN0/J+avkAD3yA4yq+Er9pUCeEVnthUNiB1ms
SRMlc3wMbIr1YBxmw6x4AwMp7Z3oFzAViFZ4g395eAz/0Q8Vhnh27dFrsDTi3Pc6/Un4TgVMrKA3
fCu0RNyV0gfp3rYdmPzzQ48ud6FxxHSvryDRaXYeUDTudVAP10xV/fr7Thq2/01L9V0sI7Wa5jQt
d8Y2Ah3i1NX+cqx3W84bdEwNJ4tPnU1CGXaaqRt/w5HPyjJ0b5EYY51sa5GqvpmAKPMt3eqi47VF
MnLPkJbcv7EQlXRW6oMQumX/P/eKFjPeTB8Zyc7cW9tNSCILBYCTq8uz9aG4PloEmemh/3tMFKOJ
6rW8LHqGAJqRS97jIN9Ahnbztorr/WqUmnGXOM0V4eX/scZPyuKvQbNBGU2PfIjw4qNqg9ZaZptM
jzyBecy1J0sMhRsR66R/p5uYZA6vFj2JLMLko8lw286mKdjhfrd6eyaMiCOetuYYm6uziFbKgUQ3
JrNdHc4EKPjzipdGtPf07YOun34tJIcOXtrMAXi8qCdz+Mau8Oxt07kqje1WHXO+SOXki5UJC5AS
IfusjMWqdPCiK4x45+IVkwTtmkqXn4yzsMqBL+fOZDOh/evWUYXNTl7rZDLytYINGsscvH6j4B+y
RtVABYQt19G14Qr0QDarwOHzV6TugwPCtgoCAcWlUgBbJbgEeRgzY5WVuubBFtTtErlPyw90jy+f
9IKKQObTG0W72konub/Zt9c62xoABkuTiowvUKidWbzZuD4CDdoauS4iizyWJ/guANL5Y4faTjEd
evNU1NmFIokw2tAgjnpcLNBwUAu+JRhBIpK7wRYr6J4F6LgvHsecr8a3bfRjnE/WVB1kFRXcEaOn
eYLRlgJDNSxcYhf6fA9Ni5RSM6s91NsUPDVavLCUDRHXdX1dJUyFx81Kz2WGUmltmwjyQeJc1i9j
mb5Mx7SYcPeV+9HFfUD6ZLSOaDre+KFG+3CU3Ls0e/F0sYO4CPoK5VkYx5XPWekw65kEjlbidhuY
l4lBdGK+7i1r89lNLPsJ3WZbJGDF11ruCcw3ZqdLD7L5TAxIVg9zUpqsdHZsTd/wluX5JcYcSYhH
C0Zx5GQIkxX8NfJqULKL+OWL6fFv5BXwib7XFcNS54Iytl9UsV4jOUEBXx9PmqMXqzhGC+GYVX69
AxPSAZ3BOTbvWIdYQNyESmWPU3gvCeFcRkT/NWNysqVeZztaGoJldoSbH0ZqenwlJ9HxDigCqoLO
DuR7c8acAGiNsJz9DBNfyPUueiy0tPl+F4ukmgU7RiRhUHSiCkmBrGucuGC/a99qvnJIcbq2oEbe
VvJe1r2+HOIy5PjAxqhTNNKEPi7xgmXsP2iV2QxInL92fln7jdBah/dMoUvYredg9ZcxuzdTZXq7
Z0khEDlfouio3QF4kAkhz6+Jo3BOPvKoeJ2of/yyXRojQEz6UkzCbIobx1MbGQJsR/PDvHWGcr4f
kSsN0aNzw1BiSgDI7FQt8QsCOhpecC8knBzKJk5H7QSFiZ7WsrHeB2h6JPvcc1IOLWFjCIhaDsnq
KiGC0ejA8cBBSs+DlY1AmO1AI6665Z9OsS9WdqeAIWAvRR9uZRuevTTYLryi7G1nhhpXWs7lDglP
Y+/W04z/RMknL8vCBwmicR5mRGsZUORTi7AOomy8dRc8g+ySX7ORWXx7YCr0P6B9400u75v0FsNv
3SysPuxVhhZJGx3JtZqYYDrEMS5qT1UVD6g0s7J0xyF8H4U/x63Tefj3qxAZHUow2z7HPKe12E0P
UWSYs4J6A8OG97zC2Nf6QXzIoYHc0/8Fz2qo/DmjxzlFzau0YMKlZv2h1a2j6w+bNjHbyeNh327i
JmXtXyoIRT3JIaJtmDG+ft/obIJ5SeOERQ+kKga84gV11yhWM7VmBFH+y1oEQN5rNdjZKsauwxaD
i9RDAZZq/53Cea2zVj+OdMYqQYTbcqEbBQ==
`pragma protect end_protected
