`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aoFxfKHiMqSEyUbvCihRZtljKPeS7PlgEHRrO33hnvctLgzxZRIHs2pewYRVwar0
OZf77E71UOdSL2Rhhu/zvy2Je+A/yw1mPy+NNJoSbHHZogLZrnS/xfTKrtu0gWdw
2kOSIC+7MpbKsYsB+zUT/XxQCqCGupkQPszZEvpwhBA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 50080)
xMhvFmy4DoqcN+2thjIeN9emrv/KwNFzendds7Y0N/cIdUhHWcSWSRsEK/jpvGiZ
HD2axPPKtFpXyeHRP49lV6i1eSVaBucdY+TuF5Jf81NryJa5fvRRfi3MfBUtUzD4
Od8h6HgusqbEaa9PvqhjIaaKwuRtYRbrzd9zxaCWWIMgF3CIWKioyxpTx03Q2u90
8sswg7+Cql7yA/2s/FIEaeLOjyEH/aGgbZhaxaOLOHibHAmOjQLCBqC9NR+M015v
i4P0Ziw4Wk6N0BJNspnVQ5o1An2hEoS4hHhudPpTyaMlcN6sfRfViXH4cT2PYm1A
nfmM2ot/yxQ3ELXiFoev17rhHAfVBjUdURumsavhnQQGI9ZBvpz2pkQczYgaKyuE
oGcc/MwOqVoEI9irPgkICcpob0BOf3Y/6ECay8KrU6MNLRH5SnSGpT0ILCXEfsRj
tXmU6x32ETOLZdICig1Kj2zkKWNfeikgbgOTDFxeoyNanI0tYZAxN5uzCiN+iUyA
peTX6q2jZb9JaGk35JYScUU0zPWcdJ79B7yaUQp346P+2rxI/eM+coxKKSF4qWNy
IABREpA19YNyc+mQf23L3u3SRg1Xv4Hj9/xMRjmvPKabKgKA1hvlXaUqX0lzXWL/
H8R4tT41sG/aEC7INaU7IJEhJWn7QIgFosxtaLPG+3JxoQrxv4R+Ztu0/tD46+Bz
qVsEjfxaHIDW9H5Ki89Sc4CdzjtcXOGMHDjOY9dsHr2z3Cd7ZLUGwgO2xpfamjQ7
d/0PWmrg9zcy1rqwpDuCGCxLger56B5HIFq13nRi/IQeOuBOixDO6KY+gIV7CGWr
KBTL37MM/0UzeTNXKL+bwthaFj5u0/YNeXwattmzlMIxj2TD9Agpx7kbYhrKJGTI
exSdpe/y+wUgDfpkmwjKrVtQ19+ERKTaa6fm0E4xi62b6+tA7AqjiZ+aj3+Aixbq
41DHieGe8xVUmSzYenjnTPZkXXzLAIOMYjXod188vj4Cqpp96KuXPQyqYP6kJWOH
rjLtSYfU81dXqDc+JBmptf8GdJ8KL8R1AF3s32WaVCAuW6VIkLz10DjuLK+ALhUa
olYPWwtepSWlIQH6YsaQWJaZMsdcgIW0G8/IOVLshfQ3yahtnu2tN27FCvOd0SEm
X18MW7wiJRmdGMW+RnwvHVtlzGAcJem8HadSkW01DbJwwTCUcHN5CFXZnwAvHdQC
1yewROgC6SY+722vKCgaltd3hilJQjkoq73zvxvXAtslVvUqCaDzCixb0bDzWI1D
e9gihRp8azZoya+brq6cPqYPaUtToIEMKRcbhludKdiUkIM7MbXZsKisUJvJQsNd
f8ZLRrvZG/mtr3vpg+LBCiRoRotqKTh5L89w2poFgfPxb2PIsZLiBe4Gs9S0/tC5
6XYMzROSNj+XryzpwmMktBE0IPYUT/hJoJT9D9QC7Ab6qDWMa0no8ZKFn+KSZwr0
IY+ojs+JSKi9l8A84E250UW8T3WzYGcEv07KNqg98QCCDYl5cWo9FxkxmrZAVvUB
FgJnSS/FocWHicI5RIfIAIisaPII8pp7M20qzsmQBrwVmzgk8i+LE1/5mMpDG4zA
6gSmfZyYGOZsMi9MhSXp0hwiANGfIPd1NvYk9U1Apm67qfR1LB8NWMDYJl27BwLk
j74ws39dfYX1PJONO4vRM6oLm7AXvi9/ny6xCSUdR+imRhuAzEz93dQKU07sIKxR
kCqbEC9LiGUvmenMOBiciMb/qf7FgWqRiRxspKqVy6dx9ZOy+RH7pJrSYlURE71f
vFi3USgXSYO9yx2NkvjfW1nuH71FXVXKepDfIAQfpy6PPTJgTIDJDlsz50lvkD6v
QPoT6beYyq4tmg+8AiAwBpXbREQFecJkxHPf8moKUNDUqRBN8Xr8yssiyLJG9KzP
wFM7NHyIJ5wsI1rYdG7DkU1UPjJtJmdr1uhbmUNgCcPfQnngiuxzzXdobjFmH040
WSMJvEYsvSflMmRDuoIs7/OuLhE9SEsJKElZ9vy8aM1tnka0Zy3zvP8Xm5jvrI18
Y1UbbUcjOI/u76k9IP54NDwfkOnaMW1W1IIlYeRPQiT5i7HQ73puzBJsUkOC5G0s
fAbBmiRxLrcGZo4TIwH6dpiUw19TuFpufFTi00g3juOcs2jlXYK5WNGdKP1i/zgr
XJBxECBOXGWJZqFVbCGlEBsMon2aB7bd1oQUcLytv4qU798n/34dcwuIr7lHzJ4y
l/UfavngolenU/uFuEsSERca2MtIolcXdAZ1nJYk6Kv4DsiN6flqCOX15VlXc2AO
+sawOATRzr6WI+ZMsjRREaA6z/uozjao6QwbIFp9xxOJPqiXemYTJvA/RDN8vvML
V3q+rvJxntVtA7iUxbG/uQXbp4RG9wKo/I9yHobqwDfS/nxGXQtB/9zXuM1fpIUY
713UvHLatfuq740+kupfJoTFzL8stD2EOXSmBDpkW70/OxRwuxLZwSdD4bngirXT
cjeKcUmcmK9XyYbKl/OWKkreeg0/bKPUx+FJy7Hl5bbB0lCjTSGoGkHBzRArmjv9
q/7j0dECVRwMJ0OJL3iFHiXkhFMQw8oG+J0ywymup2ZqEcbv3AX8ZT7niHAR2r8v
PPRH4o3EGKE2e2wZotDWxt1zpYqKm8ZWJ9Yl6mfSiGrSlFgl2wT5RkC3Qn3RhIA/
UCFI2K6g1n8aXphLdTwOLxDRpSsRE48GRiX7N2PAD9QjwNnsmk9hHNpm740BZWEP
RD6zQ4iMjT52O17mkNQSkI2CkCykemK5IDGpEFfkN43edLPHO03j2zhLeyQqp44T
u4LAeO06yejrBUC7Hw7NsNENexu9bexgGOCWFWrw5HgZgiyt72Dz8/fzo5snz7QH
NX+aqo2tM15RQysEUGaDCmfdg9QT0xNlodzoU+Yk9k6dQKnVjczS96SZR/WCTsed
WN0a3YQKe5fvjVXMvrhmIvP3WJVmeG3J6/yi2nXLZYdgvsWaUxtgMrEc+yzVyp2G
mncODGjdOqUAlBPvyq//Pl4CX2o1yKiPOGrP9PiYDaWC9kcZ656jpl6yn+JI5QfF
CsNsoJuDqhpGBreGswLS+nxoRblpTjgjKcXgWmTTzO/4oYV9faHYSG5ySzD2UT10
ZcjbfnlaBRwpT2TXkCiq2DwRCytoFhGzRdgvXlLzd/iwowTtMQIofh/g84sDWRvv
dd7jkzO2mUF5Amt1A4Z9DJrl/igcBtBeVBDLRsyS30B9jDRy+HhqXy2zVWHn14JI
nmI1xLOwON27STnHBjU6kUflRHUh7LqpHQDave+7la1+3X8LdQ0NQgpTofkmMern
xo1VNkU+A1AFiORRBjtVNYs7U5bnuoN4JP2BLrJIGm39d/nGtJB/KlCLbl0UkMsu
GBXGxCM6AnLAgsVsryoBNFh3uzKa52k0E3XTh9sbOJ4inSbseFI2Unamp+REz0we
sX7kwZTCFxnEFyn1mthk+XETijP2sTKOLvo2nL3a8HJ7CEVwQzk5pd5dDhTGxdys
g1NVtz0YtRezuoGsBKXQ1at/7BI8jqXYQ36mF07jBBFJhXmcNWjGtoVZeG2opcSw
0MAoypuvTbYQbwLGsUweZDHNvfHch7taNbKAkSoD7rWxIZ5MW2du21DqfB9PpUC2
Pm0GWMqBt2c7YodDvoWtuZolrNXrw89XvTKcAkWvqaajBhp0Rn8iasDY1dFSoUIp
JHOda8C4yFdvtJrlmXB8S2ImkRnyqopp5BPydRc1xnJoz9EaYlV6BpTbg9Ib9zKa
IpLCDWO6uMe0tz3Xrlpeldh88hy7XeHxlv/PJr33Hsf9BHWI78gKiDavDIvF9z5n
nc8UnnqoGaGaEW8aOyFlp5u4i68AcH+UKU1SY0ZEHsIBGo6Uq3p1yY1VNIASMu4h
Apwa3gOuC8msrBMVGwl9YZZASReopN5l2xEnmlHrfGPS7KXpOCy40B1MvCGiYmLs
2FjjcCa/U6BDFb/FMomc8VaLZM+UJZEte2k2L7/Yvr1VZEPM1tyYXQkec8a3hNJa
OZalMX/K6kIMd4GhimxCJEIPlu9T04itBT1w6jixuUkOf7e2y8ycj3KhCy4KiVBP
nXLxslfgYQEzH8mDR6okQGucQZeBW4k3gkgc2uHP+6X7e9KzMM8/O//Bk84a/CF0
tjoornHpONWyFQHkMzbojDREau+CHGUEOepF7efYebQ18omA6M+JIYo1zIos4jkC
TZ4oI2O4pToknudpfvdUMIOowMHd7kj1YQ5Ei8bHXPueI6QWQ6PjTqZerg2Fanvk
XWucLcSIr/CqL08hX+F3D90Jg5/y7vK7bK1Rrp8scyARm6k6ZCJphsyTTIvmT635
18PRoidCcfsj4iyrTGP6QYY2gpPJyeojTErWFr359LGUd88uqiqTTTzFrwOD0Fin
+DvpZRxOjHzYrrd3405iNN5T8GjFBvBsfhBsrQ+b6otqc0uhAU8WTw9zxiP5IpMh
R52a55Izf3vo4LWkGlPsUYJJ5sGpeB2WE2/wN6elxBj69bnoRro2lu/87V79LCzV
19pkjf3ZlJP+sHSngolh9DXv4ACuHdNR0t3L0NyvF0iRpwE2RlkDjEOFb5xIk1gi
P71Qq45UFFPstdKqnoPPfR7Y5gjO8HF1xVtNN5vuaofWGXjFMAQPUOSABUPOXX5d
8MqarqLpcEy99LzNUFEPEKWcMqv3xezJboIT8AOJB2/UV41e3tVD2mzebIhjxL4k
zOHEssibo+ZoSJ0t7uOr6VNmc0Som1sfEwKlfxY4Tl4UeX+n8PnULvWUFwK2SvWZ
ZJllIt5oXOa/FXxFCRXFKGdKe1qRii54pVv1nV6ibijaOl4n1b7U7Dked4c9U2Xy
y6ToS57R8sGIGtQYd4ora/RSc/ESpM5rLzgYewBM/9KGpkaGCyHJxadot2iyWjn6
SCtQNV7ZsrwV4t3fvKJIJaTZDOm8Lq5y71ffKn0x5HH0O1LHHkOi0PEd73uHNAqW
yjy0R7vl18g1zNsekiu3AC953wcPzFkF2ZX0s8GIbUwDOjGZTbSM2t2rxQ9KupcW
NvTU3IMVNlu9tz/9RT4D6TEDXOAWPb/k5i6gdmy55xkRrHt43AFlGMa+9ezERpqc
MLdydkV0hvhw+5Y70aMprtzoi3LCyN1sW4EobehVzO8ixMCn/H27mMnBjLV6MrZ3
tX3ddox2lTesVnUrGGSvkZUJag/P9QYNT+ieFObKO83frkMoaEfWj+iK++BVSAsF
VDX5VhQLdSS1OXNnaNBLrEk7YXZj2S7gy3+fhg++l897k5g+2AeAs7hkWLbUFSKQ
u0oKtdpyxS/oxsbA276JTkx7PyrK23TqgXRRbxhprgv2/OZDoledO9obUEbflZlz
Rzm+nkfW5Lxygafhgn6srWnxFoHMxrBRWn9t6AzMdQXSvo0TuHRYzKFJQa6A+1Ly
5lZ4hX0t5n2tbuqhKxO9T+B6e+Nd5L+80YPtsSXlFDMqjLBazlpVHfO6Fz4UM9hN
JTPFrfD0DTUbpK2Giuf1p1Yi4uLDkTdk9yJI0bJnUpd4MNdh8Xsx51OKPnSG1VQ1
Y3YzOivNBHlevBN5hzKKRALhqS/t2MQlULLAp5pkjGyIoQ/vlfgkm/Yl7YOxiTjZ
6W1AF26BKbBOwo2HgxZpGOH9USyyssSs5su9Jg1l9VBqIdCrDkw1MOa7H6U0JjG5
Pbr03nczZaI0nr5j2Fo3RaRaSaYgC6hJ5PYDHpRGXJ3XD/I/Wh0ncYY54q2VgtNw
RcDr0ybg4guzbDt+ETed2jL4KE9wkAZwu7Q7/p/AvDbp4PlqoJBguZ6C93Aht4dJ
K696s/ICz8k3yKjKhqklhH0Psmcbfy7xkROhKZZ+kSuU5bWdIlen/Aq4p/coWtgt
96B1cmimtkc/t6z4JdR6F2qQBuB3QLgzeLE+BtB9bV+fnnlBa/7Wdw1H9teLHitB
bh/qBv/Owpz3PsEyeBAtlhUu9eTBSKYNrSpQG7RufubDK+1A4UEPEwo6Jq7OYaj/
eL5ga9UQl+umsOles5wk9KiQhWvTJ/+wEtFrpbQYFaWNcKEqesChgW6RCMQlRMsC
VUT3q1xwtnQIkKslw6NRH/TiOMnk/J4S7OGy5yGAdoVqaTw/2qg4sjOohMe2Fc70
PN+VStR68GX8AyJGoVMYrAZ5qne5H3nGGp4grmrqJD8COm9qtgfMdH5DpTVR5x2X
9GPSXAPHwPOwYZi8Cz2q1sQxN71/IwqC2CdGv+yjkivN6bo4Olmnr2ClcpujYxwW
wtVC1MpxdOBG0HH0mweBn15MdX5oIchptMmLGuLcU468jJQB1CP5KxzcHih019wv
mJyznd2Tsnh91oEYozjYEMDFDXzuaXRJLEyXb82hjEm6jWSY5qnEVcgAhUkgooy9
+5uOVywd3RHVLpwy6UY2dqi0wvxjQyf6GsAw7awhfDs/qyPXwZRiNM4cgVBJLMt1
jCPbPwIM1y0bnBJUclfBmQT9RBdonQUugVSX8Ze+fIkJHEe0HpOM7yxg4V92HNzu
/iqRNB3ZOH9ta4ZLt2hiq+DNv5LmSYEo76vPyH6plfhEuwVc0UIqWY7bKt4Z7WPL
8aJ9Om2U1gYdHzs1ll/Tgkk7sw08xbPDLkdERStMWx3793jrGpd0NpcUq1xw7nHn
a0f2Ij3fl+NjpTOULfgm4eLyjTK6gJny7FNca1BEB7+zNHTQcxNDgb2Y5q2KgWT8
mXG8WnLIwb74N3iMl4TntXVT3FSwI++mb+53+VsPCCjS37+S8vlouCDf67bUyD4M
JFhNRZCjNUf0gtJp3WmYwNQURYHJCOJRt1YYk3v2U26+0lMkuhDV25FJB1rhlTLu
/fv5/fx/ueo0OrHhd6pLcOipj5F56KJdoiu4KQLv8TBiB+wsXZFB7KGXNZTAtOwO
i0KQeOk4qX9StZNUXZkBe+vWc6IjnGnk5rHwNNJ1QYvd+4mScKNBQyuJvZ7LjjiP
u4UXFFDpJt3JYjxylOdWvmdhrLxDVmRkxJS4yUAO6fscVVe6mEQffp8tOK3woqNt
UGxaLP6XjGSWI8YvnBhUVh3FJsHOryYwevxC560Bz9I+iWDv8OpcddAITLCT9Ua2
0WK4F3KhNhSy68cfjQRE3BSPgWiVQJyFW/LW3IQXty8/0+/lEg39CTlrgoxLihl8
SaUsDffkCpnLUs1ULkVfVL8T+TwTOj3Rn82W9/yX2NTJdDW9sYdiRPxoJ7BI5Qdd
zQciEWiTRP4/GLPI3PLeT1HrvsRU7MmLOgt9+7NhNztOkwWgqfqZQtiO917cJR+c
ZosYBJNCNzEZifwBJeiX6TBEgP1T5fiGnnm2fd7D/zFIB7ra8pUEB0P5rOJUAlyI
z0+hYlUtUIvXLisP86FRmSMfdIbxvfUJYArUgrCRgCxjwGzCKt+HMicPhk7DkYsJ
kyOt+nf80P5SrnXExJP3b6ZUpkvMQ7Too8aQNMmnyh8XPRfWp/IjzTqjdb4VKePo
YS/DqECcd/C5Uq6hhPm87oDbaqF8G83bEkcpFnIvTcvxPHxBvJr0SyK8QM8JqchU
AxxZnHjNAWyu0kDXmJW9HUFrED/gE4LOv0t0wAqFberH1mK3Yli4wPj4fYDgsCn8
NIyJp1GDTnY/CgqdkAVbHiKN60/XQ/26/MlprpbvIWibtCGazkQEjt/SpWEipQ8J
QR49+++E/QcYNAv3s5GXxov9p/Han7tggwZBnwuz068T3MKzn12w6nUODIlEzE5f
+eCc/bg1owJVvAo1Nws9kjSHwEODs/OSnxG+MQc21+ytWvpbO9M4QlxGMhOZN4OT
xc29rvOqngeEqqLZlAq5PqSO569369mCGUANhLAE1DUBR0BZrRWA8DiZfzSIRMsr
a6/aXBpJWDmaI5zEqR9N5LiYq89452KVFXc1C2YMcpTOaHLRq792nnwTxcFirtod
Sbq4oB0to64GU+B4XKKi+LEE4ZivLUCNnIeUoMOWRhj+k/hUnxXzQDtV+nfsdq+V
Bh2WI2Box2EX77SXgLPv2zUc9VVa1eASePVgZsiL+dsUEdyyJAPmfqJAHLXls4Ws
Bpu/qGsBprRNmr3R2bfs1FfXhlJ6T9ZtMFZQaxTlP8msqXFbsnA9SgNqGeu8TSt8
LwIEnCOD0P7nCr3A79Yym4eiQM6f5qUoQXCG0EBomndXeysGz8kBBdSRnqwEV3CF
9drARyXDmc0UkQz+nRoRSBUUTRSN3+zGdO5Rv+c9AsnSG1zN7wraYiXShF3vPhmE
llzGxh7ehRjM2EvIxw3D+dqSbOp1nPcxcOr2P9OWxVa1ssmqIzjR2QuKdnXTGEA1
wMWDG4Dkh31/Ng/ZUVJVoR3EXl9Dh5foCw6jKOBYfjfsxCEAEoiku/iaU33ySVoB
qCwPWKOrOs5DLnaqV4XmH2IXsB+PFn/ZFqks5cfY24ofFZ/tY6swTfqlVKIEtKl0
/M0au6KBtv5ZeJhzAd10tG8onndfOSg254cKqR8PzuCLGuGLbn9jQudfDTITP9+A
8peotdicgu3PM6C1h7hRQlPwQnBApvs7e29Pbzn3FV/JrbQ0NjhI/ncOgxPrM0Eu
niMnCxGoi73AQ6xbTV6FRoE/4AeAdyn7UfHGog+ICHqL5FDabJooJef0yeZWFScL
t+6YpethQru+1XyP80h3Yi7CGF0Husf4o6oi1d6xFHD9MHs4ged5Innqi5mh6/Fw
obh7/8d2jhcdUJJMZqZCAmLchUCrdrEolSzTb9ToaCM/sRDXwiZg/sMtpbbNrAna
J33+cdk39k6EotrQzWt/iHdgKa+p+v6tJYKhyv+6d1ZHVLE2/Co+ey+psvL7AAgk
VaGtZEnfgIQD/aSr1BB2RFHTZARpnT6EILEzlXwAuszkylPQx2a84eS62oc7YWYd
sLfLVef9x6hpVrFDUf/IHNahDXx4nDjpKa72MIDnNAMNkmMEqX2x7in6XJf5lhgY
8vDiNsk1S8XVOKubv+Z3qEQFbXCN9JJfqV7SVMXI/4rMn+iFVnILT05S974H9nEx
Pjuo1ocBEYwR6VY1ixu3iJdBHdX4FVswteIbwZVZazfSaMVPP51DGKR//KHXsQ5U
TpPrurzGEntOqEuTU0QpNlxVd6xlwisQdvo5dycbylQ4PKefeMgICCJYG8RnDe41
NQRQoJnHLpcg/k9BMGw0NaR4qw/utBktQHP5LwzQQzHFLTtAYSdMROBMfik8Ik8e
b7AhKiqgq3R8uzVo3+HpJr1NPLkSx4L5arfte0QIWvUIdikahnFHvuDdepJIklsw
Laa8oBI7CShQ3bkXOIQyT1Rihm7lFKOVUgmZnEKjzQYgac4h5V0VwFM8rA4yn/o8
m5MZ7jPwcjyWJXDNAePjuR3Y58SZeSOqvDW+XuYK3p+2WO+JhpmVAMSM5A6XRraU
LrQ6lV3XiT6OSnm/7uKE/TbOcBKJ82JHXkplcSSkSjNl3t3ho2si8oS0KXxHgVDm
Hrz44Kof+SQXgp2Y9jF9zzhZLS0bwOJOxMMeufGuLs+uE2UkxVn+41JJfYv9v3CD
1iGuri5JbrLVC1zghsHN9zsJgY4bQdHhMnquQ1l95qe+6f4Owt0wpkve8T4N5ubD
6nk7aFYuAjswyLhA2RdT+tfMRygvfsos1hNeMz0HUL4eE6HKMzlcg63aXBC8UVqs
/vpt/PMe6PKYGUFRLQr748hGpHWZ0L9+NVyuZ6ZyK9V2spzDtuPPs5G+G8tzHmfj
tyCzWvL23FQ76KyPJi35XTSWCPjAdGB7ebLT5St8Wrdm7YnZ/96atHC995Z8Bbvd
MJe6F44y7mZDwmBwu2ALXJ859TOEN6qgSvfVCmTRyJp39OLCZxk+cdQfd/7TUCmi
HkNi+Lk4EUEqn/3uVNWw2wm0sIKRRWCueErN2iJuvKI1/Aq/gbMZZjduXfU6vQWq
rkxsSXmocq7uILg9lVVdhsKwY9nYhnTU3K/yOAt32JfkCIUI6rIiMoo9pXyq/90s
R93LivmLjP1JhL2P5FuGAThbuZqUkz6ZtQDk8ccprgzUnh5KQkqMQKTK6nC65tk7
pvxGaqHdu+rOxXHhT3DXTgs+qBsgI7enFnDQOJuxx1u4lqF7kzU1nsMx1bAclB5z
kSI6rOj9t5TMlNKfr5jmeujGh8O/aeLkmJipZzWZ4s2L139EEEAWiK/HLLE/lxLG
RfwLVebCzI9jmi0HxQxdlkFnEh3MgHtPQzckXdqiPQOh5pq6OrsIWcXE0MSJxnQh
fYt11hN2ERggyQDciT7h6waC/pdBMiwawRLVa6fvtG60Kh934XHYiXGRWUklrfjk
lOZWsK0dUu6iCWml8jHt7qFfJM9MO81EVm2aeFLoxpUfeE6Ah46LbbceY3HpDEQR
SFfvv9WdjZZc5eHgLYe04RP040LrsU7LiddbP72UaoEB9k0DMgDX6BAK7la2KIEI
mr/e8ppZQbhsRptuaMn2q7W8jeaQKqUjLChtLBgTu8cc9PuFReB9fadY/4XGlB9A
0Lfnn7rAHzPpmJo2u9mLAgQPKB+6aRVmO9ogeWxBYxH29c2M9pJh/FkyBe7le/Kt
G4x8D4zXZH8T3ox8YU8MnBdRBvIVBpGnRPJEmiiMEqLC/SdUJEqvYr36R3rvMe+s
Y/2V6hFrt+9JcbJY3aWZeXZ+IAVKbD6Bs9AidrsL74kRECZOIijp5+AT+qxlY4En
4YOOK1F8e1pGKUrbOs1/ff0UirSUzRvi+DRAe/acMi3+vL577XYWR768XbhOjC9/
W/TjD6Xi/zuzKq7tCSg6SU2H7M6QlzxWqh7JV6bx2Rfuc8bJjESoS3LuCHy/XDUt
CZqYFBhrFvuU8T5Cg565rJv0duxVFmwOrvA7A8MiGpIItz7usIUpVitxMq2JytOt
Oak57vtW/76r4SDZqT6wSeIRsXOMJmNMOPlV8Uops/tzjHcQkQ30q3bYGsM1Wrnk
AFmrV++dsu/NCpvyX1be8Y9l5y56+PPBVmLO0OuIVqkUIPHAvKjvxi7mdP2ukFxF
uqgmZs8VwswY02WeSGkuQt5YYXRfYksxu7Zbjhj3qLLqLntbnpZYeeL+JBt+n8QW
ZMORkxP+ZCDSZqV1kOdVzf/8sKRh24zsFg90B6BCiiO9pov0wmT/RmD1sIiJzErM
gWv1yKg58G7/Q9g02fNYnosaMiFdm1FbLHw9OA/+Cla39E9EI6l1C6iX/ANP7w/k
elXLAyJmDP6inqDAqCeQT/RuEN8xJf7ffG7u3G5Qw1Dp94V/sqvJ8k4m2OV5UFTi
lx67/G5mcVM1tBoEQ5J8biD1WXvyHcMaH/V61faJFzxfIvVQaplwblM1R99g02oh
9QDCpNd72RFv42zYg/afBzFtrT5MNfziW7cotr5pQG+7YGoNDnutxFxHQAMnIEP4
J1TRwyFJ3W/2TlAZVP5v0grLsDLmGJCx+QjLGSzyLNnYx5Q9WxXhnt8IxDLPSg2d
7Df9obEUL91VKq+DIAcE/PkwPFG4sOa2HphKAe8HZCeztIT0U3N2cwIP3b3Z9E6l
fcNfQumRrQ5f4HJgCms0OoAGEd3t7qqhZYPI16s73DQQgnjYeL7fwV0b597TbngT
UXQrdELRKjW86P3W6K1FtiMZuqRfOqB4aZxkhUkH0nBvcrOQnJNC2dlTkybBjjSI
6PvfX7PLUQeoY7iOdV0nnKJzeJ6hn11+OLmzZb2KRi2nSfbfTMG/vgaAHc/HieBf
Phn0k6jfsZt70eKlxEmwGr6tO/Gi5TkE/OYaKeANwAma2Tp/IlZNYUiseWOp304q
O+u2Wht7HNwDO5mJt4Y/lJNiivS/qvqdwQcTLzxV0OwVFUUedZ4Env/HfVBLA3OB
pfcBn+LMghJSdP/11EX+L2UtpXED1ZoCgN/PTprLZqFnHzIIxwAdPLEwnETAEKlZ
G6jGKvrIBjImtkbEGkhodj7N/cXn7RqVM0kVFttHbWK6hreVhSgOE145xpY+PpVd
9aiYXcvsTXijheChMMLA0yF32M6OhMA5UiAM2TiPcNoU2srA/fpdkHOT21xpjPNX
NpGt3EGo3Dvp6J09Xs90dcFVMFYgSJUyzxIPJnOZkATguUGp/7qeNCyhdvX5qSoO
5w/bdvkHVhlL4jQqvZjJ/LQYx8tiAuVOUm96DB0mtZPuxEAD9J7a719rOm1PCWb1
2acqLT+yIB/yQL5yvRwSicHHmkTbib9ehO0LtblWTmhJ1DOap/ABfCd552p00ndu
NUJv9KE1tPobhlCB5tM+nUSQp7bfaCPvcWQErQWkcWCt7UwQ6TKJVKv1vl//TBVk
SfDHf27JPxj6KFCsfYSHVrvlgyw6dybj3OeiMhkzLgzg3MwduxgG50fSfRDf+AkB
JOrjVv969cZPd4vOsPzOgOA4sYtD5H4rDqouNxifzP5gId9Rz96ZzjUa7n4xpZTG
3/BX/hzb1iWfxnK38tKX0ur8a0+D3YkuSJOKRth018a9z67hGLFZGWxnXE6gGbci
OhUsir5f5Mou+fUeuoxGRdHkfXmBcrvZx0JfLRC2DbPOM1Bftr0JKRMdlKne1zLe
WDEtxGi083eivqZs769DEndZxYo+ZUBd4Mkqxou32Tz4uPRwQbw1TQz+H5NtgITY
Wo0HI0ys1KqEOeTZU8pSUZogo15AutaqqjAJSX3GSfahEh3e5ju7rL8CsHpg0fNA
rF6FeCCJq8WnV05LeXI6ts8UokLzNBVCYgvh+HdFhp5vnKIoFN1ZvEwE4gNc1I54
Zye6O2Ed/lhWmxUwd/30gMzIWtX9BbiBF/FIriTNEHc/mglRLl2hoLxgxoPZXppB
HnasRY5KXVNf9L2EAHdzeeiu1JsugsuQ3GsqX+pHU+bpIRoK18XG7Hl9FClrK3Kr
GUDqH6iXGE+5RXkUgbBnIQPDnYoR2Oap1fTZnyLQAmCpjSV4l2rgrQZci1PHKHyN
5VgDn82VRBTQKWbh0zN4ckzCuuW1oQnpV8LykO2onf7KW8qHm+cA4QHnmnJHwPFm
ofW4hnGXsiVk7RZMAUnGTcp2UVoZ1qIvHRE/2kxK4DoTqoCuPmoZi02YxWla3cmv
91tyzoNRqWZMUEargk/rAqKc7hrNa8+e+JVlHFKTsmuirAO5aUBAjChBOShAilqS
nySq+EAQrLzkaRFytOJtX7z9qlQwrd0lEo+Ls4oi9mAm/D4ycK7s1gwgt2jEXQl8
g3lX1/LQx0NjXoI+U27oD/wIyKnyzxvjF+WpfSpA5ML8HGXTC7STAUcxAHhCS95q
mMmARS8GhRpsXagMUdLyMvp7hKmkeQU1462PqLprnH9q+Xa45gLFarh3frqgQkjQ
Lzj9fXKUG3GLBruDncxz/IrOoxpOgFvoWEIgb4AuObolnGNNygu/JPzQ5artcs8Z
1ClMJSNGSdPFFk3BINj+LLXRTNS77b/3rB49Ym1U66kND3LktV0TfAICD/Z2jdLO
6SqSs+IfJcofMkJlThJphZ1s7UcKPMcAF/5Z3RbLRSbs/x5qjaMxYj0yBGb/1KR0
RZyL99yRRHdDq29hvo+YUKs6rtpvS9adZQ8fgHirLU7lnvi6OwZyCiisOGsrwbJ2
wxbyS04fRzMWjeI6h7ytit0OYJrln/FNLrMF4haL755bQm8qgLVTU2JIUm3OIjFH
nO76BOx4jysmF48yrkofNOdIgD8RmUBaazW8Fw/Pl2+4LZcl2vbkLd+UgH03DRtH
gxoazEARlgFZCXFOaiQcKFlLqdJO9h6Q5CT70djb/I/lf8VOabdKPMW5oFpW68jy
5KMGVGzT/Ksx1psN0B+Xue/I0vGiqn4C4Xr47uD6Cl/vlhukdTJDPHvEgPxPOi25
6+waMcynGRwW3N0tO+JeKIdQpAXg1XgfwKuDHy/Xk99DNcBlQvskKgk2UuM8cMh5
vS/C0z5dTw3yuODEK/hXYMSN2YR3/pSFJtaPdpSjFYTCT8h9AJNInjVAVsrhuE/R
uqBpLklxzDtCHOzGIwZGzUU7pg3bNW/aowIKTkxw/61POA+8XAo1TfWUbACCd67F
KPn0mOuMuhZOvCgWb1CaM3nst4lpinLsK4yS06fbCpATyD1Kx7AB854DYgFgrwDc
6a7zpxDZhE9SuZKY85iTNJtPezGoQB/zrcp4O9H4Z5MR0ckYmUcYmWrOb1hDp6Kv
3HsxCpc9y1plgy3p9HEtei3CwHoHiJPPZyQhdO/cGLU9abF+kKu3VD7dklEQ5MBN
/OmZnAAApPSz3qwgf99zED4ZB1SqSQx9/M0gDkuT/hk2+d7KmsDJ2Thmr5QzxZw+
9dAloFU+HQhhB2rfzPDZXZNqvgshRo38o34gJGs9ECjDoQEA1b/ZfPh9kJSjXHtD
aHHTaElS7u2pUwKYMXaMs7/qBUKo/YR95Czt907Sy/Y0vm3mV3IKuw2HyQh0V37Y
wbONyllZgY4ftepWxaB52y5EFjt+x9R9M9vRcEwDAg0vBoXoSeeAGDpeq60W7zc/
OmzgrV+Ye5bYm0RzaxC5s1m5BiZO7iI2oIjbGK+YggKos61atYXEL3IveMd00Ui/
elyCGN0QqR8JDik9qQ5qL5UKKMsdMBN1o6GyWq3RRpAcUsSlgIArHmmE0Skg7wnB
WgMzqwmlhStxiu5TvhAfSS9ruoABDortP82ySQHLGBLnF9msPTnubhxnDgoZQjDB
t0Qt8R9zRrA60R9OS3W+4scvN3JD6ID604jetAj8/FHeQ+kSpDkRelP2aKS+Q4FE
IWIPSlZESGdTVHEN2bhA0Pf+xeQDkTavwRLK7VRCrAfAVbYEtSlRLxI0Mg5lySfO
duQdFNmBvyQfEFvSzVv308cP3mml9K2dOIdhKhSt3lTnZmSkYrXw5wk4fi8flT81
p3GtCsP52VvOAVXykwMW81WmKBcSjTYfKc2xY0M8+dLRRFXLfgyIfTx3RGcw+oM/
n+zJTa86cov41EbLtmn6FYLvA8VeL0qrtanQ+lzufQlJoCwtLI9O4AIp4W/a3D0I
VmR4pbnAetOGptvuJ6UAgX2I/PeI1vEwV7kw0qxRm+VBR9WXrLaj/dTTIhZnfX5g
feJQ4sAP/iDLruZYvLXMX+eUVipJXcIGOSOfimESc8I2PuvWK5TrtqYTeI872MyG
7g3rw/yYpI/p0ExXS5Qy7iE8h6l/ij/q8iHkYVZhLZImkbPY+OdQAYZlffI6BHde
EXt6aeW8pXuupf6wTn3MH8tLHFA8k9wMLGlAKa/TFXtS+ifjUHn/ZtaSTHhD49QH
l20B/SZsAjqCygCwO22Ylj7bF/2UObauYczWKWy+oKXT6kbU1oWnSmvOrjI5zQZI
kx3/P0YdoPR+QDLtE7y9BFgSEdAlcITA2cVvPFVZFdY7cM46kw8f+rh7Q1uuOUd+
ei6JLOTW/IXTZZzkYVEEKoiPtL6ylPZGq2nuQsYvxvw8d5gxcYPfUcItN6Yq78/H
lc2ZxyHJ5V7T8xywd2BDxJvqzJM5cLEB4rpWbuTdC3jTnB8ipkD5RkCQ9cpGh/9b
53G1sNXUmzPdkj2JfOkY8g74Z9mdOm9ETb0MfZX7L06URRhjFdIfmIazvyzcOylC
PR/AI0hm4d1qxuxLYbyB4GRw1U8GvkIZt7p/mp2Izbe+k8y9t6+GU6zPvAaNKQaO
evEhGzkDUaS1Rc4pihYcEianY8MWTOmTh5SdeujUjf874Hp6QXfXWTG9F+aGTpTH
GRCdKrJGqXUJ3cqJ6I92QmlOmBeGzj/UbCj006K7dJsRoqQUMX7+rpP5dhaPe2ci
OCH3y9WeLIEnJn65zMFT4pXdMyWagq+jaTOXSKvlBOI6tPpClMzrpUtaCZDJ9vOl
eu2lEkc46bCsxSGdGkHAPR8eB0HkFF+bn0sb6NtvhjaMgcQ68aWhlTopXzv8WJRi
USi5C52q+Lw+ZaOEMPZZLjC47RZOkneFSfTmll+JXD6fM/0+3p8wW6lw6z0VbXNz
V9azGOaDEckC71GCmMiZw37avluTWCKfMGcmHdTN9dR1Djxph6IXaL9XPDov9Ttz
CSUWdX/PZq5yZwIs3cnU+Mrfm6f4GSzrfQETEyyGw1057pi0UL8ImRnYUB7gLtfC
r3+Bf5cuI/70NOSMtqQ2rxYYbeYLgxXhghcPyvaZH2og6y6VnwwzYUfDJyEJWyYQ
54JuKuZa1Tzr7PzFJq11wF9KfPBOHgxsMVJjlbtedLxwkUb69YBZBu0bxvkQVMls
v4zdy7+12XCADlAu4XmzJLaudeyJBAtJ35HFfWup53mfBNUKy9t2Et6JR2OD4oaC
BvmU+FmmA5c74guQWxcbgQ5n/y0rPYvN0UrmfkLgktyzI0pcQUDN5ZBG96J6ye5B
PqZRIdr5EXVuEqoID6Kwym9t2UJQkr18q/7tVa6CpfkdJBBg1g/DYuvF5uZFXNgc
SmRhGQwVhpeHuXnMO7erSx13YkiQyXjTJ4Ky9aeDwBj9hqvDnxptLeCr64wOarH7
/mlruicp4lZLqHRfHoLeprzhKPyA4jyV9FIRWsKL24EoBYX2v8v+ztv4Z5lbMhoK
AUdoS0KtTKlC9h7B6XmFpMyhRSXSjilP477kXDBRp1FhnW+bv+hM20M2RYPPcgOV
3eUa/bj91uVIahZh3rl6A1UYH8fJyCIEb4YngNY6WsjE2IagcV8axPlvwudT7TxW
69mvgKh7F9exizlcpeCzlUzCXhSu0CTIu53oeKzMZ3Z6B1PaYCgijeBe7OHVUwGD
QXtTGdbrR4jzoll8sSzqyPY7qtqy6QH57GPmbyr9A/ueiQ2EfRdXHDdtW/ZqNFMv
EgiPS5WygLOoFAFdE0P1iAJ+P7hjzwmGJ0XU7Ym0mu9mkQL2RIBcaZLKjjnp7odB
BtkRRoKKRKnaBjWCyS8B2ZXfGHPE9jQlt5Ux7PdEfdjZ/K6BzHpEanH/XNxalm9S
IUyE6SfZzc/a3upvnTMiz4dpsfr1E2FZAGjtP/HqP1faiv/k8S/3MjzSjPEyZmSk
ZzwJlua6nJFhd0tL1JcxtqlI4/hNSRMhYdktqRFEZuQn9c06d1KWlINp5w++12i8
YjU14xCADWABdAzpfe1RT7GYC8xEAROWdgzNC7lbJwo0yluDC+67IoUozymRng4t
WIohVL82aabvCaMc0QL//dSXWkwk3xV+i+wbynDpXWLobDIPvM2flBTY4hgzeFpm
TgY+ze9SURSJpL4jb0JQt10/MllVLYof8RdW6s2yxvW/2T3zEzzbICro9szDjOOH
9CTha2kAj/aWe0GuyKKIXtAKuB4D5J9zLTqqjUfwknIyZTJrJfB1ItGRUFZgVium
PmSIG/XdE2Rtu9boss1SPrPNpg10VuzeRnSh26uSAG6FCjqdml0W0+JgBqZpvZ3z
p2TJx5FoKtG0ay0opb9EWVDmGANsNuI5khtAmc4FW1QZmVqKqCgsKxAut8H1B3sk
zDaqJY+d5KgXggnZhDXQ2lM7+MhNwqjXT6ElTegacQiZblJTBnIaCGH5MTcOqLks
+7IYUeXxsKQg84Pa+W+F3aMK4LsgrwEM5LzvjuTLI8DLq+ipoU8cj/7lOGhw9QRs
EZrES7sRDQ9tTYneh1f6ikHhiDSD479PRfpAKRU80L1+lCq/LIrfQrw7ex0CDI8/
3t/V0t6foBTinE9tSro680dbXbF9sht/5WcppOeJDZsq/XYfP6ep8Ki9utOsFK9D
wcrzehO+stYVFDJwJtRIKuynnqhlb1UGyLzCSciuhYFo7LhUBMZkivX+oAGuGN5n
ylq2LlxO2QFlhASyX4MviJPXazlVJDnFp7F1jcRAAeGagB/cYLcOk3nHoqlZA3r9
vqrBnXDh1OtSFsp2vwYIloIoxk2mvsSt2pvGkllr4SCSTZWOLRqJXvfVfVZHrxT1
YNaV4mr+z3/DnYit7kdYdhW4aXileoTVxbbwc8x53e5U+ChlE1AxtHwjrgn/I6lT
Tc1OLqChxNzC4zAFdUEQu2lwfgNgOjchQUSIenTwRum1B5owdFqfDMqFQUCbwV04
qo4JL/d0qkf8mPLlkC8NiXRfjOCxfjfLR7r2isac5FO4bGlQ3+9xik1zy6JW3vNT
7pguwPILBzkQ9ZvY/zqoUtezdBy1xmH812vruMgx839e7H/KneesbgB3lNZMN4L+
FoN2Kob1C2An1q6jie0v3tm3qcMJbfjYHDoHlbJLvdF/WD3pQWBfiqSCgNwqE63s
6DSqts9gDwUHPLP19VgARVATTJ7iaNSNa09kTt2dlfAZabVU9vhvKpIpBy45Vlh6
WCS+KinNdYYbmAAlY2oWICDcvEPo+6Bu93gQFZX6r02v7T7A2EfSmiQ7X3bYQrb6
sHzt28tFwju1GX3tIvc8FIkgS2i62txXUcFAxuwHMJZ2GrSbG4TqJM5MT1ANQVtc
1IaQbhVSPwCWq+dbkbNMNlks3Aro941NT8e39nOcECjP1ViIDUD+YdcsTEMD4ZXt
CfybCtDW1+DqYrWrXJM+aLafQq9odHtc+wIJl4igtAZwDXBxTDjUxDFNd3tfNEwy
tCS+rzsP2xZ0wmK/k2QfdCdSSm8VfyR8VGy7IWJn31wDWJEsINTv6xpDXVVVlMSA
7L9/sAv/wo0PQB0D2AXfG/d0MwE/6Yz3hOGXU2r1wTLzZEh7CzSFeqgarL+gnI/9
qJm83bPAHdjdpXr4HcnrfH5YiFxAhfSOhcjq1beo7WjHchTVIcDvF+hq+GYmnQTF
pc4nyWRLYGwGCf1VvAo5y6P/liFCgM1rzl5AiE/IziZR8QGBNRoQoBZSVmiJGa04
bGWxmImPZzCZfBDXGsEItXkERlIVIyZmCN4z5oJMGc+F+2m3tdSUgCRDotS28itO
YJBtvFNzR+3riJK+gY7owkJD8bOfVG7/Z/0+kui4C/Y//dZN8cTxExQIF/mPrJAN
8C9X9Egm8EtHK+RDMpWZD+Aup8Ya1tIANvEntV/EZI+ROZp2mAcPDTeWMKbzQOND
PGSBl6q+EaDqGqreFHr9UtGEYFvgrFLepWi2duuuXIjxZOmbNI/HO3LPfDG7DPzQ
SrOJM4hPimMhJRMRV2zGsXw1PAqwsaz405tnNhrEIZK2XlcYIqqxNO1PSbseeL0+
PexAfbewqfauUX1jkepdLZrpyu7T8U1cclgjbXvKxCJgcL/9p6ONmd3kAZnD8tst
ORp32yu4qj0UAz334PFvrdm7EtxvVHvohwrTpjt42xtgc4OPh5hk1sA4JJ5sGYBk
fezcON0Hk0iUyd9rUNB0VuYjkoXaw5NBCPiZw7cRP0gblsnnTHQ/PFS+bE6mAeQn
XxJLorVHpe7BsFImQNC42LO3C6JbOyktNCTfl3tZczZiaqGlEARPJaE0fV7FPgr9
m9F/teo0W0E+/KTSqEMeFXe20WFjqyoYFeCXHfS6IbM/wxB9cfQOum9qrweUZVwl
cCG2ku/JWZgZntjI9XNVIM+haBHaH3WcV/o2iJx+lZaDxaDxfrLRLH+rlD0S6eXn
aAEyWOSSUWZcz/CFXDjZA4ozyW9cc1w+sWa7G991FFvtelpF823/gp/G1PG7nlCb
F1773ff9Baqy+5CzIvKhKJ4Z/FLhA6c+H30oJcDgZ7M/lk5yqhEbVl1vI1Ty/XdS
zkUMCXe/IIZ413tRwFr1yIz/24gKBBWZOA3dmy62T0CIZV44E8JTx1f2l7zw9DIL
IrDF0Mn6brhyvVULn6gKeAap1Z9FDTSAM4BalT+mKB0mZ1p2cp7qh4SB/6FLb8CA
fTnUBcphZBOsyDnO7hTN3wiwVEhCc0MiGXcBLShdH2273oc5NyOMRHp4Yqrcy0HA
TFNG56fe+9txej186LrVZcl9OB4EmhtWAJd0aF4qw56NumhQ4VPSEr7g/xA/eWvE
CJ/jC/n0FpjNCPOj9TaJtys+DyjUrpNGGCQRTTAGv/+ImNu30J1iNLvSHsm5cxhS
ZQ3qPb6Lp0kDa28+HUJxr0FlApdpXshGfycygACJ5JOsLrIJAJuterKVE75rTPED
93U3f23/fcOvJbZvwcDPLXU6cTfyTuEdzaXUR4s8IiJvyIc4wDt4EI+MMJUVN+Qe
5NGHy+mTajC4k6qMwh/5fYFm4P75NMz5YSHCEUZET7fAtapWd/aGu+rNaSmieFKJ
v4h3p+pdE58d39XEWUeA7foCapBqJpRR2sKrpaiz656LtJKTnAvDqM6WwterWCu8
s12eLHkBu+QzEdHjZ2vnIEiInKZWWLfmGC0VHDDli2HwSVHzFjfu01s4cAOEnAgh
nOV7vG6iRV85FHV4fbNg6QjPr7tc0JTsEeaKcr4EQzuHwLTbf83T2ScYewKyTQWL
d/VhrnIrLcGLC/MzRpofG8yQbhHDfewWeBgdDdR9sGAAOZu+Za80FFjHfS+HJkUu
2wdYvfBJ5WCbWKoJBVcdEUlihyJpg2FRg7I/WonEH7WaZgGb0m9ypTZZoVO/nkVP
/Fz2EVqcGc1r5g1YQtRe71DbP+6j0yvdB35kvm8fjaaGADyy7eOxST2QL1QRzqn7
tZhPM4P34VgAiYdwNChD/nzjPEaUF97qKS+P1SIZfoL03ZG6euZL2/m7yOgbFBPD
+ZsmVklZ16U8e/toowOm3NjajrKKiMDj7bG+ELrJFGvsPAiMfdmB8Db1J49iwbn4
5LrIDP97HdaX4RP8zp/Og19d/0cQgJKpb8KEQ9M0vcMSG7xlJvvBjEYTqvn2v7H9
qFeMw3t4olgC3XFqmOfidvDVYx03AZnCg9OwbbLBtWORfr3ItqplG8fqxXvnzaw7
mxu4gwoiB2qqfr667DBlRYnSfihwfBvZ0jtROeuOvBaFKFDxJK3cc0PqSC++Uda+
p//u5TDDd7Y/hip+LGLgIDV5gbge3K6I6AkT8+yZFQ7pNKOXBHrjb+efvsB0axYv
z68pZxx1jgQV+ERJZdyq2/UkYGBCzmxgZuw9lCNTMqNR1+fBUls5nxiCK4uK459/
SJlWkVeywyNnAA9SOacS+mUDIaEsOE+e1drNwOOho5CzsxPh5QGItcjK6VBOPl/B
Io+tnmfzlk8X9XdIN91xrZPT89yVomlyNVu1ynQc0s77Ksq/ffpw3Arl3EPvkRmw
cTDxNtDS1uJaFnyjCTLUfLry5piMk2HSmwFIoq25kXKtvLr4mxuVEA01NdWyQAkA
pdlRY3PAPCGpGVbRL0JrSmyAdfv95JSZ+4PNUR7NmknMtjjeG4FQhhH9v5LqeG0u
QbxwzWNzQa1O0N68xNoirI1smWvtAM6NC+NCz+1uleXRhGOaes03wAzhx1qVbS+T
yLFUU1pLUWNc6WoTFwKBtMsWcYbw89i9otkWph2YsHiz8eIPaBGhDp3Alth1CrKe
iEd9slbD4lV72QgmkgsEZ9F193BzNYIjuhRkD/r5oywi9Aq6V7a/nrnuYxr8hsLD
8smbFa5g69KJqtHR+l/6GSqaTUpyq9UKOyD7op/MIp2Zg7PIVdZ7Qh07sxb33XqV
Qg73atVfZZdxH0CtGU7QyT5L5IS/JI27zjr4GLTz7CWgEopLIcrV4LBXrKGa6BIz
H25m1pO7OvOqK6f3K4G3Hdm+0/3+LfHp5X0WCLUDLxDgEncBUicOcSRAG2il9MwO
+gpzrddFuQD3JPeoFLns7PTk5ugdD/cCgFInKUNlb64UG1cw//JM/1SxwwsKOWAA
+z6QCNYNTc70LgzJtTjUF/QgRtvkyy5M5oc5r19QnRKe6eBf2eq42GmlxH6kNZj8
Jlki1B08DyeuzIouyOeCsWcsMN32g8AOfHNI7YuVLeh21qesBW4KsXNrnnbRrtCR
C5kPcbFGcObvTR9V7ccJdNSqHKDrykTwMDOljinWcOQL81XdkQJgaKBe1LUmM0Nf
su7/K+ysoHQSCEpiQILLnJUIxbe7fWmFk2aE9m/E1LseppR+LK4E6458QiiinsqJ
RbI1Rs7uWKgc9nAO20Kprx6Pse/eZibl+jSVZ+O197nGk3rkXB/FV+YWyHNNNbLO
8KbaAuMnMZNVc44dUEvJCXDFkXOQnL6BUb771d8g5a1LMLnU+IL1DBuqcH3H6Vp0
r5RgEltaOR5n3NkWJRwCOZwYWSbQ3DAPyrNj0ZsBdPVYYOE6UHnjw8dtQX4v4tHo
f70xU+o/nPs7vYhTnIu3XfHgGVMhyCTfjmYXfz+K//Kgqm0+msfd1VTNR9mdQAgD
aryGgKxqWvRcPJw8h86Ig0Jr9FhgWonbql1xF4QMe2dlvB8jXXCR+N38l5Xcd0b2
tdAwaRn90BXN0dYDAd1iJprR61RGCVAK2A0ctupqAA/iSvc3zLOvAbjBS6A3rF6q
jzJQSujQrOL1tnvoV8rSSs58/YsZ5ZvJ5jhaFbvhgaseCSZdj25GnrYY3HzAMzER
PH5ZT+6Ajr6kfHy71+dbbWsR+YYmyE//J59/BhpR4z4qUdWx/hr8usPuO1DjSy5K
BJqjA5xaqXd+BGqSnFbtD7xH8VqBn1MpkqBjHRAWzIQTNC73muVsZKmza6+AYEL1
sKTt98/lMD2u76vLr8O+dJFmCg7qKWXrSz4Aa+EhVYqUwMdb2trWIaFggAni2nVU
LnaJDTZERHrsRYnFE6/iHQ6f9c93AZetb24FE1Mh8qfoGy1Wb/pYNUmjHb9Qn5th
iCMcivFR/86+6kkl+FiMmmxF+so0tBZVTG8RYgYgqdKNcb/Ksr/UOTA0UX3aC5Po
99/hh8j0nScaX3au4kHS3TJuMZIh9lAu1g1nOFnfx3V4lRDgZW4zzxZWISEaRR++
vk6fFWuhynxU7y7NCTzSYsjMM4xZixKxbSDW+U6f7O1+fE4YPBflQGZL4B5esF1J
a8VJYcLWXejTfw1U9xdRbkGg5qCNC5hD6H2YACOctg3VUdfdk30RQT9bC1KDbDHU
bSH5qd7JCZhjYjprRq5sEUpP8eMy2iAz7zaV4r/Prj49g3kHiJlGypgjJk91ooKv
cIaXsVa2EwgoBqX54m7+BECbC37W28yZPod+3bLEpdM4IaRKSsSlydiEY+hTc091
7hZwDMvCKa4qzUsVID97fWvlsYV2s4jzqwO/bde8ckMT4gnI5MiRD7/HPVnuuTUW
oa/EIUGYzn2wWSe37K7ySkZkblsvcCOb4bMyv0RZiXCp5VM69Qt4BsiNQU1yohwS
/3fA30/WTaqyuMFDYcbwtFedCYxC28h199d87fsxXDM5Novvl4gqmJBwBA3Y+9fZ
ff59gfOKZ/aR0TRD9AlYi3E0UVBQiKkAq7Je/U8EjGeBZQ/7dCz5CmcSNvLeZLy8
rpqKyco7oyKM29rU2JGX8u2G8gFJ1MgxUaVVw9/3peHsPaEMzSQ+Msfj7x7nwtIH
FjUbkDckpsEXebtCPfFl/gIlS4Jy7IFqTFDrR/aB6f7pv8PJDaQlsevRCW1K3RId
dKCeh2EsP8veIhCgFL+WEc9esXu46gsdiHM4wq+hGLTGRXkRZTNM0MK5JGT7TiqU
IkK4KkviDWILNF4FB2awZtTl0S+rbaSuFihS6KjbrlJrSaLF3WGNf/W4XTegnwd8
C8daGYUQGwtebcDphOGZegRQMgohjmcxGAk5FXSorFWCLy3n3apEhBTGpvCqCd7F
L/45AAEvy8gIouRzZ9sJ+b6svo2/hd4Zvx5V8K635s6TNFeCnQt6+jeudw3qZ+oH
4qhSOxr1fl8DEiHBm4ls/S2iTzkfGwxwoY2JlLiTxHhV4E/tdClO20OxiM2Rh/Tw
j1Rk+mzP2D68W9GM8BJLsl7grE2SQCT61LdW8gY7j6zsSk55dzxI32VH3SqHrDsu
sY5m+8E5YCN3KtGn9eou8EwupTMZha90yeP29WCTH5eTWx7RPackyLTCXPPOA3jP
9l3vk3PPfCKnGjFtExyAYOqoeqDguRfSaeiccJOO2WzFZfioKMVej2VW/wDDJdDp
k3aeBhBtg9AF/aZjnvsbWkNdx4UQqRDaGGWEMgs0LdEW0yPKXoBEm5T6BolR61Ct
JQV15etjYFlsDSQKJ+Dohz/RfBmCvdsM/PmRDZ681g97eNdccDtgs97dEHaMRMpk
l/sqzB4wnRUoTPAr7DVDIk584Uq2ABz3aSHc/8BVV8i3J9yajVa4/SRibBSHKsPf
e7TN4VatvUxtK3kHsQLVLjFguwoeIe0Z7T+zk+0qfCW3FrbczoSkb60XRkrDV1+x
cfA2bHdF8zkdLgH59srHldx1zLl77gaoMgDNyfuRKUtxFm+TZQOoJ6G7dpfnXkem
EIDNB+p12JAMRcnAdvoS1Y0B8xtUx92J+l1pDVMcXHATBOLUEXQidJkX9G5QNT3Q
Ikc478PViPhorIBzCq6fBTts7ZBtDMYfjLxLH1OrfQC9hLbKmIFwx0jyRZyQAh9B
xyC+dfPLlJPtGlGF97SFBz4boJz6Rx/+wsNMYrP9rpq+phNt7Tkb7WzFMqSv3CL7
UjtjK772mLIY4Fh5fC5kqqY+pzPWp3gJ9uRzLarOD0xw/6Do/KLT2RymcLwAj18Z
+QrC0GVlb4/o4F41828zub5ZSLnY8vMWXzTdLFQfHaWqyIIfGKaHgsTw3mhgJ3WV
OBIwrYlhXnkhitjZ8W3uOlPc0RxcwEEiQZcdk0DIIU+biNzShE+NPktF6dIdSLNP
P2MBLS1qT2BE4azHubF5u/YNPPdtBG95RIWujFuWtv1VPMgQaOfLnUONh+R43R0L
LOtENiFccP70YUXGLiCOD5cxhbtxfCkN58pkIk1cK72dJc62LiiikONgfX5UF2DS
YL1kDSG7DaHAgo3NZ7vCfkc1YgjUP7gVqtsLd6rSew5QY0PXSbhwYH9jmZWIYxuI
Pj/olrlKYTR6Z68aCvKI5/sgW4k/8G5Kjk3B9sRy8ut2KbWgSaI/XEhV7lHhOOua
ADoArO9IQUOobRCkH0AqjezsIe9rysbugD4MtreOXZjroF9n3FO4Y2KYhSfMCplX
bZkk80M4X3SisxVmhpk4DNTvuoHcdwgA7MhACFN25Y7tkn/nxaSDC5SVwkCMBSpi
QvT3jhWCGsZBZqLAlbyUsGIh8Q6bwUZBWrW7S+wYjDsxU/32aeyMtTWU7G1iLj6n
eT67DaO7OsvlupUozi0EZi7OxqSn8x0sW+saCfTrmBZmsHmE6F29iZJqR3jcl8ZP
rMZbBcaw2UUjYuwF+AEW4n2xHCLdoIaaptULrB+joskTmEk62Ux6bBC6qb3vq3BG
zXuPceTsM9cpESPKYSzxojwWbyG0nNrRaL6snRGvY+aMyQefms3k+CrSsIlC/bxz
MCM4AO3f3Cxy2FV6wBBoQ2brV76iNMLaZAdThEjx4qhGzHhc67xvZAfHJ8V3fw8d
XFgtTfifl79HcfiLrj/ggQTULqSsx+69wMIRxM0NdGyOPkBTsNXbfmIxjzNKG8MZ
q79RlleqMHXOdVCpdD+59/5+jBCMUbywXfqP3Yw/KPlq4i0cMbmXfjOE5kx77X/8
os5umg9qAJ5XL5mBEp26clmMFe/3Fy/Fulgg4td29LXAzt6yX5sHqVuHmJSVuBGN
wczeqMn77g9pfZSvt/skqf1qJmOLo1XRbD7DMnGGgpcxDpD0d69Hbe7PTMu0J6IE
gfc1WSeqa7qHglxfwMw052bYhp3B83kxxDdm6MUKR/az8sYvFZFWzY6A7/xw1H/Q
GI14MAzIIejNmFue7dz9MHXduK8a6S8C/HJ198TnACq86kWZR4NkgKQ/ArFVf60u
tDyMywyczeafgnNjXcldW7PtvNqimuTjPhO7ipT323eXx8y2kU1IM1Ju2F/6afTT
ONGI6WJ0h1RYegf2VQBrYjYYIBM6xopH/Ze46xo0w5uOUyXfv7y+WroTWU8BXXEE
PRbCRPHlgzkNWS2Bu4vZI/Ixfb5MzLuCaxS1NzyjiZeCg+4zVfE3e1mGcccw9kJZ
5mGm68gG2TYs0Fszt4kyL667wJXKar20x02PQ0X2sCmtzx0vakmwWVSbMuoPabBv
SB3CHHApMpVXYBwyt4qxZjvm+3qPgEDJbyKl+RXX1x2wehBVKfshimNMO/XAyrUL
13OQHUXIISKNWPFl0QTu5ulz25/y0CSQatjXBIhN0fgGDbWl06C0W5dSfT4wR+Y4
Y4YAoNI3C1PyNK468oF95+TkQYen53FV19uak3X/RxhbL9M5i0T53H9+6xcJUQpL
ix+XF/NKp/M+/Q4jyCD0Cl1whih0HoMQ9nHs4502arhRfeS6wleTRPeZorBknBPu
ZbsQWqGkyCBr2wjZjyfv9+TWUC+oH9iUNMapfv0he2pulbopeOPnLJIwweHhWk42
9KRRPqkjiBMSmBN51bYezLTnm+aAF0wiIh7yXkYdPgJrF6PUpPlCR7R3STgF7T5O
zMRm/baEfh7zzT7yS8f5mct6tQ/4y0oDeFSv62J98Sk5Ny/9oFaXLRIi29aTXcYF
gc4zUd88EONwmtvKq6imNXvzWXRIF9Nd4DQ4hxGrcJk5ZkflXjM7soi95jDlNNFg
XnF1jR8lHeueWwt4Rjd2W16D3wy3wiY2Hqy9ojLpDB4NtraxU1ywBs+o0meyczTq
Hg1Ilii7i/qkt9ZQBnmEmDrSGhTEEHfJlp6Kf4i2SM7oHAS2HM5FUXSVYO0/0mfn
BlFb9hz0fFPRBMWAmmg2tun1crOBgiuczYehFIj0X4wn/4DCR5P0+ms4768B1XEh
uQxa790asj/sIyUoL/GxE96mGW8E7f9UBPCC9LAu6uJrHWwi7zdtDnueOhvH9Wi1
yId5nTd47wOJGvZN9SV3ExUiJlw/01nG6FV+Hd7I6KnsItoJdg+fnjCeoluS0Vfe
qJxgRRTpIjikif0iCLUczJ2k3/J1JZ1tdgK1fGLxd96H8XUYDkMHGq1Qx/bXTOXB
S0+hVSyP+k52THdyfn9XLNzj0XhX72/xCi0ScjIptfXmGOoon0YgeOPcVaTG8T/z
dGwV0DZ6lm94XSy7l4XhqTEGoQIHun4UoCeibvr4xJ0S+PrrcEAcGMmjAzJ8jFcb
BNQEKrWMjipvmaUpno/U8cxNZpEiU3qxhjNqUEPayNqsiVx2PlIhpCurypwX+9zG
hECXIdAlVlo7ble7Cop3LF1J0Ww4DVP1lvhLxB1XPRMXrp1skoyLOXwqDPWUY3Uh
cytnPzfHTNe+2md61jy5DqSBxwr3vhqBjKC7cCUIhJewbKPJfXu/u51pVxhYczRu
USq50F5jVRkLdwR7W/odySw/ueVXGkK7To+OLElbXu1gtG977mmhHk5jKT/WLZxn
KKkcUFu7aatrxaobjvsx0R/Lc1jD2fxoCYDUYixVqUJE/zLmBoF+/dFa3s9dx1W8
IcPi+xnHMgSAdWP0HEntW0Vnej8mW3qC2OWSsKUQXkmFsNns+qK/UpndO1TCL7vc
Rtz9eU+FQjOcU5RHbUQvtP9Xj4jhjMsn+Zd0aXokqM6wQoxNzpQFMIZnY73qU/Yd
O/yDg4sNczclcBgWoPIv2tshQM/sKdaYddv6OUjMeTNDxqROIFqJPYRk7Tps/dMT
IzziDImsEETXmRR4L1mEm01N00Ca4lsGCciBr+95d1dC885givW5wrWYhP8MOPrI
3QS4c+iv4LSbvSCQS/5yh7ml0PhBI6KvKmReZ+Rj20anKAJ9fuQKbU/LxKKZ1Qr/
1ymsbXVR9ImoZPLusqi4yLwrEprv7LztVJuMJpHKMDCDoBNTeMsaTxEiAVPlsIG7
t6gUJt1VltX9mFhhCCySu7+AJO/wTjO8iLmtRft+/l0SNoSyn2i5JF+qJbVIFQ48
Dsd+hyOsnK0rDN1UmWwqE23ZpgJMk+lJOyAqckLvpzw3mpW6+tyXZl9UMhQCoHMX
l3/Vu8jUxp7TXxhY01vOaU8F+DtXHA4pUUFlzLembFzoaTTyeusDSEddj1xEwalm
tFULQ0q1wjx/u0I20jvtWKT551ZmyScffiKrE/T7y3r89m0TTU5CGT4WjkkReO+4
/VDPthDiLwvIhoQewSbPU4lQ46CBHYsXWt6ne/1ckC1muCY+v81cJaLiC5wjkyHT
4R4Ql7C3cqTJyrLipxdFU0hjKjC6bzBu80yDWtfUb17TNuXWO5vBGT9efw0XkPPK
0j4Cw1CUd91KAN8+NwePHy0pgUXqjLKI0aJrFqzCM3Y3k/TFJK+gM45keSimCLHT
QGTZc8MddZMqWvQ4IOzVuMgeXMdyC6kQPCseb19uhdxU4QqQGC6FJ/QnxWM2Jh85
cMGSWQo+jkZvyBkwcU0BYG9OC4DY9vZJ5hP/GA0bSZo5J8WL3V6QocWp8G4Kw7DZ
4TQX2rxbFCoyi8adVylROGarZneIvrebOtQh7HPeVaXu8YEi7HYu0Psk+NSmpa+f
t7IvY9WRhkd8eFT+OIVbkZPbydgMw7yPCtPyWjoORQ+tZHDCCMa5GCZF4ln/d6bX
sK8qyN79kQm6j6B8kN2MMJhfyM+ritAIGI4kKWEJVZz8NNFJvQqFn7QtqjLtfeSi
9wxiY/mJDH3qOt8evkdB9zrNHvkSWiIvEpYONfhYMpgWyTbXlUKyZYSsKQJGQlKj
7LkvLNZTy2gpCi+qbGZHQ71USGnP3r4LJzVNo2ztf1X/RHWHpHVuuv0ZtQoErr5o
rhSRKRy+EoorkHFIgg0NpXJReYAFK2XOrj6JO5CnNiWwfABVjpjQprv4YNOjl7bz
IoZ0mA4vuqixibyKsm2kuRlEWQv0S+q9CTCplRjytqHaA1+cIO3vpqTPkRYGQ4Bk
GZt95LVO6zE4oPqZmuDxfqh4Jhquz27T+PPkGf437paszCo4uvxldEpGrBXdYfeB
J7q4JOIMS4kNKlAt/tHmBh3C/Rw3+/bn8b47AoeDAffVETS5Xr9Gqq0jJ0GNZ8us
XRctwSBSx5VytzCUuGvCYz79fjivQjHTbgvlNGsTAE9wHD0l2mu97hwnZnc4a3Hc
FEZcD+VI9Mt3R6f5rWLxOEM4Hx26u0nS+RtmUOJFArCLFShtMNM3ctXshRgonLo4
w/BvTFLh8ZbBgiVlie1gdBXr0WJY9iioIXv4JxcWFrsO2JKdEytkTvNWW84/NDbV
Mi3LrWeKzFkwGEZwQrVag35dhAUlv7B7cBA1pQ43riuH2CMCUSbLDBNltN7icSuA
wk/y5W+0hloYCO/hpPbLx663+EVtvTYVeetykAshiTh7UpQBoicTnXKTR8SzcRNu
UYEViZMyOwWLswhNMQS4qc52dqf3IbHjktNueCLlWCrzBs27RB/tUoRePmHWMy6I
XaBSIiMFyBE8JLs495//0M2CqrGdT1FPoAzwIkxuNL5AVmrlZ5PxT8Zd2K7ms891
xHWFSA6NCjIqcnBmrCUo3WthCmYJ4TGbSOfw8qFE2tdsd+HouKZHfE5242aM/0IF
pIPbfIV4mwnRO6unNMXj3yzdWCHZfgsxlVJmrOrZ93FCoIXHYxmtmRvd9BnV8Dma
fYgIQej3JNaMArW2HLMO67jlJXg+C2nRG7jerS94SzR0kC+DY/3Al5QfxBRqPODe
YTEcUHpj++fELaSwWMXIIcr6uFfhIJmbD1wuXBfwC6D9nTTvhBDOkCrGqOc4sVe2
SFLNI+Wk4k3XuaqkpWukzc1BR/aRwv1VtiHFysBBUxRVh9u9WUmFJj+C86o3L9XW
oyOdatevNd8baH0tfnvshjFy6O1uVBVspM8GxfHgMSMk/12wsRBjYW2uAvCoGjmB
1Ous7CxtESQczvcLf/Gg2bw3AFKmUhWwm6P9CrjTIeLPSP67UmaVDp4gj+f3jxKQ
gCA7llmyhiBQJN6auFIs4jq4MV+8tajtd8ZEEE8SBrF9dnJJkzVrr8cDT0PDSi2n
5v/Envx1JHwrMytj3vM2joNOCV+Zfd5zmbOzuALAIKVuWy6xooZl634XA/2EmTx4
GgZEkSqFj7lM0zkYwrxA8ndNXMGu0yf8x06+HUhhVRXcIPH15iJX0fBDreBBvfz+
WY9INLDmWkuwhILBYGrSCeCyocOizT8mX9quJp6MSrilqTu76txvRotCfxePxxSG
xVZNPYW9KSnjaaAHyapwGlC8fkvytTn1k4NoUqDoQJtYP0n5OxnTE5rb9wmyhGTK
AGTq3Twfe/QerofN+EjiBXjBjzB6sNFrkkED6MzPhBF4PZl8aXARBsoFlzupyqI3
glP8+cp6gGAw/RmhbnaxcJuKF4XPbSXzvDydSETk14xjiDlQbCIRIKkQ46vanofs
ZMbYDrQedokgYpgyHZajp4yIRhOM3gkHCVv+r8y3NBaPR3nYAY4b+BJwOwBOrdm3
C3hvhV1BQYed3OCq2p6iSb0Sv3ZF4UJkMhxKcZVqdTPd8e8R8Vx7jIP0stm4xDgV
UKAF0C9tevSl2V9Ccbw0KM3/o+JIURl5nMlmCp59p610tESU7BsCAnLuDntePNEp
n3fRfG4DKNM06P86R8c7VSMlu/DzmS1VIqSBigmB1btVmEZc4jZbR631EuhevYMT
tOrp8Vuic+uYCRAKcrcTLXpnMWve1VoNRjRbJLYYSq5F9ECdZIA1u9W7FyMoTKG/
IW5vv8rVh/MIwxxrFewrMGHYLwSR2xeBzlYd0/Ma4PMv1SMisibHsj8yb9TZWpC8
ZjaAYyt3AEiXwVeFQ9UwxZDMX5Qmq/OAYSIZsw3l2aKkk3ftkhMOIiEdrsgqp/2e
FGK6IPOyC+KJtGwB2d6cZXokpEwJkaww36ZLiUcv8+CO0eiUDx1w4aASpKsaSy2V
hpIWQgDwiHGGs656S5qtPK6ujE+RIEcJa5zYfEBcTbeE+v718JHACzMOjdODCtO8
r8GwqUAZdJkKZhNVwkN4X0QCMVtQzPphM7Nx60Aiftl0XciuYXWOIjiYwYU4cj/2
9LISUcZEfsdI85SmrEa0JNPGnVRKEOZs2NOECzMOWGkmnse0MKhnDFY+uaxNyisl
YwJvBqZ7kcbq9AkN2DsA30xpJTwTymEYGqhm6YiyKVauv5SfXSl3z5UpKFdv6N9O
35mKD99usH1mj5pc3MZOfYOg6SO2roNQCdg9pLxlTwJYMvlMMsaLZooe5AnZ9APO
5Lt3qeS9lIDTiaKDHqYK8QqZBmbfsXDQ2M15UjQPK3rJhu6lDDBQrqKfrWFKwDeE
g4OQ3fvvrLJhVxKHUyHIYDLkuahL6O0VYodOeACMsHhCo4loM70kSQ67ac1vg2hL
bmpnc/RDiSII1cTYoifcRGbjLtj/eoQugu/qLe+zndg3RKESEOo53RjEa5PNkpl6
Z4BwDie6J+oyLFP5rYDRBa/jrOKw7aVob/GVGQrPaBw5Kw9EWXFNM5oUxF6uRYIw
vMhFxSeKkOtuxHa9DX4gJhmSgXTzky2RwQkYTyc40r6Xw5pGv0pYpKzXQnesOkKq
TZouKMaTm1RBwFd3ztUXa9mORK1ruSBPwpf5KNpnaD3hXtq4tg3QrfYuVYCXguma
LNYC+YkCXUA+Tdiz2sqbrZ86fLS8JYXkBpZ2W0LVSvWvjV251cFi4H6eBcYlGwjn
yy1SNUfUp02ZWSGdicP5hRb5bpL02OByoN1k+u8C4evPi6YifAz1WIZ7R+meZI8G
dt1Rn83hvEKtDHe+C1srUc35xDq0l/IgUn/PdkWN5+ZrgYHSP0X0bugd7B/x3h3J
ylQwdi+1lS9TuMhmCCg0HBiQX1Wfao4eKRQ6SptPDQblyuK9rs1aflDXNK0a9nnC
/EMqPjNUnVF3PpAVFUQX8f0UEintmk2zuE0YXMaFClTKX/9y1+7qBJueV1ZyCYvy
gSq3aEobFzXCk0v7Pf4E+Wq9179v3lw2Wh2FCOIqQnJaIaukImP6ZNktW1umB9rg
IK+vnvYnoQLtrk5CjpphF5a78qqkLEw8QiCcspzmfS7765s1MbsuOEmL/iqzywnS
UBelO5DQr1nftgPG2fYL0sEzHtg5LreJaco9y6fPh3wMufmEKvSdatdGxk41cIzh
OmvDl2l21aF4nN3fiiBCRDPJfBxjnJaN+smQ1A3cosudBOTf32AKLXTRk3mNYgyj
BRDpCCB4XEF23ydGGMiUcvFix9DVe/yofJLwDoU9Bu7mNduXW8ELSZGFSoyx+gLC
dlddIgcZXjass55kFm9H0CWsYZid0Lz71yHLahuQFPjQclCZ9lf5gIW2lqWum2wI
hakUnAR146G7OeUABow0p0v2x3/xxDvOVG3Xvnb/2dBiv3xpAJpgir43ha6bWKZt
kawGF410u1TJPExJg5rLkaNp0Skm+tyueVEI1RLHf/viuPezpv48PzKr0w8NUmu5
LLMY1c5kMKKERMPSn+dKMepdmQIdJB64o2OyDOfRRYxIKNRX9uw1beQn0OxjxhnT
2L2LU4Q3rT4qDDwByxcoHYNhe1XcDN4sMTleOXepsaxHiEEHx2bC2S10ZVqjp/+d
9d4ZoJcDCotkaCFwFtZbO0dhSWzPEINKotXfpyYwGK31kJjAlLD0ktXPkzmqql/z
ZrQTVV46b7Ei9dB3oj5Uwhh5xqv31kGxKiPDpjqWAz+OUCZ+BSqm6yLSd3WOX5Zj
6RN+4Ao5ukGcLk9sKCmJjRi2Ze56LcczpY/aRIfT3DmvLb3u+cE6EPu7MAjl62SQ
wT7aaj9yhstPeEjfjVvMM5teP7WLCppTgyq3xlVNzlbCiDl8q+tU7zK5gjqh84Sg
cJ1cvhQ0O7epXkaesnhlPGxFpXClSobZYPO9r8l2uR4YXpfhf0ww79QdXeNuBKTx
VjfgeALF0pd/M7ptK8yrquz2Geg4r4PNX5Jpd1/KKKhTYrRyQnAKL1pumedjLbFJ
KTrYrJiko8mHGPTBX8OUjqSHClN++0rSgDmzFkwuho7/TldPxfCRrvNl+pnOZTSL
vfs0TrGkVCYMKf58TWXDLTgDcHOTRGiDh3Ka+UJyTgtozyCPAr6xsIQJA/+41rt+
JZ9LFetXn/8utJvdDec5QnVr8h7Uet8zEVmyYAYSr/1P9R7XR9Lqbq3McBfCV0F5
wh/LRk1U9sv5MZ3bNxlEl0HeiLdi37l5V6fX1pd3jneuQo5CMf4KXg6KDEdTLgcX
FXQhyE8on7OGH39MHSy/xwPzvUETsbwOZ+jCVkALC1+0GMA6RMAmfiEyQ4376ZBR
RECDW2pIO8RxbCqNhdnF3KSSjdbdkXhJ+P/og4n0Ar57wCcYDR4ydaSB4BSYY+iu
QSfvkXyEl1tiSwk2HHMai48yyHFHEBJY+9zTbqczVVkLPrqE/nehxYVp+DI3MQFV
17LPowGnpUWf9DhGv0hKhaNJ7tFeD4Im2TZd3drSZhZ2EGgDGIdlHsAQQgE0BXpE
aNZclo54Su0KnBFQMU39kp68OkyK4t594PCCAtg+jBxfNNgWLLj9pgJkf/0yZRIn
bI0XYzmGzs9qM7WuTsPRvTfrFTqPfmR+qaauEeudHgxR3sbxrYOR6RrIQwvyIIcb
VLWNoyS0SobYDjMOCHX6eZ2TRJBHFMiG7L+GKDEuvS4qSDXiQ/ik5+lRFg2ker5A
ickWwJnr49T7Xa03TW5Fx5Fstl0MKS0BAV3qSBcoQBGoImzN2wG0B1lkqec3D6iK
pD1QzA1+RQpmNTpvsamBXfhpD14Tn636lMgIqZjfJDbCWwlMAAVeGvbF8TnSzK5D
eR2kKFKpkf4CzN9708qadMdySGI3X02yMOVL9fDdBVo1UIvbiKXjJeUsbPbnUiPa
YWThpveyBotiFPSHizZ5jYT10MiGvPa198QFOmzQ3MGLysYMhwqYpHENpnrye8VE
snvhAD4ySby9ELP1apSgXMEJ/dV9zyCrLhHUhTw1M0sN/QnHdbL2p/4oWuTQdtZG
feWyX75VDdTX1nF9jDp/2aXoS9xGOGtaO4EBoOIBAiNRxPef1UfskjvPeQUxCRLu
bVF+rZO8w+krI45cVT5FZq4nEHfloKq536AOEzeYatlFstNTZmpNR5V2NLWTBbvq
soIeHCT5L2pWiHoi9gaHEeRn59MdxVkj2lJP8HXSqeyffFHM8aHf9niF/0uDc6cd
37YnpmfpuzdFMeGbNoKHHXDXYJAJKkjE9ErDv6qeAkiorm5zeN5V8H56CIX/WQkK
uiCYNGXyTZhAePqXH0+aPmg2Rz/YscanlZfWCJwllhAacPtAwW3BYwgCl+faBc6p
J7zWTEe/5HGOnwsfeZxeDn2NK0+U4nRf0WdR4jqMngyDxJemNSAVGQgFN3K/FTI+
bpLuPjthxgiYW5BHqh7twsiLZy9ovoitsZdgT/wwKEtnA190RiGpdmM4Jhs1IO3K
PULPula6ig1+9TQGJqmklMJcr3oJwFyfOgt9TLg9nxQNiKqW3K1MHFMdL8sjUY6t
h+1y6PbsxsShX1Bpkv2lbRbN013N4QTnmOiVm3WNlAVqjBJ8DMG7Bh+MBEk2nFNg
TyUfOyBsQ20hafy3TgsCPNudbQkfBNxvwn+KQrjxS8l7ZJNjDWtDeaY+GI+Yl7OT
ROXxk6XOKAha1U3qHnPU3kCHvUoYaauiOnnpb572M5r9PXs0TZq8Lk3A4hviaH9E
dFEM4Ep+wxvYoLHR+PaAdZHKmnNgIOG3XT4kKSd7ISXK2xJs07/wGfWOkt9X/tMM
8BwpDnFkJAXTR6WRvSgcKj7rl/6ZRBxlLg7a33ExI859HNZ/M/3bOkCshcO7CM/G
N550ufynpgMfHKI0u0ao2opfOwW+HNEGyVFO2tlKKpFhee3PZ4BgtPmOAMES7YON
ATZxaLXgiDuH1rkakvMeFp2E5Th/97RF4dP93VnKxLUYWu2hiXn+rh0WxYFtz/+9
4ONWtUN6bISOC297qmoeeb+ygsVz3E6k1MOaJUR3CGFlVZnw/SLOfytbumqWAumm
+a/Yt7D2SzgHwGIw5CAO5ky3EupibE52sA6PZtYjKxUTw5PfLBzKP2q6V9GLoMzx
USlBnaN6vfPltcup46jvZXTLpjnmTru8OCLeQLQR7R+ElK8wH1N4oCYVOWA6wzdY
IZdU7sBASd3jTvkFZB3gVQ6l13RZU04oIgq00H9wXlshSaQMyT1G6g5FmiV5VXQg
bnY2gG+lqA+AZKUljm9H1yT12+BgpO3wfxcSJA6K4oO7PLpFQDm76iLrGIF0UIQR
jOOpI/OVR7gX7nqPp91EILLoKKJsHLBF13/tRq1q6+ug6DLG5O90TEEXqhAkEcqw
fkH5Sr38ekaz+xXD/1im2f0X11UXlIZJ2p6Bapr0DSvkm6wEfqxLZ5Be42f2HKjU
Gxv/6H40KYumeVaSDE6Zwe2dzPXRwvxVp80ML7njlSttIiSYgKqGbNShOFS1Jynq
4pOHJanlBIuupercRgo1ezyOpFQEL09PwJnJa1WG2dQNMMErgH4RL2FDKSyzXvfK
U9OwLhunrDH/A++idX5RIlKkPKGmtG8a3u4K6xHfIrM1wXTdnM6i25rdN9/q0jnO
LH+tJSYRqPyvPFElgqAhf9OTMMX4IJKEkHk4YYOYRrzPF8wgESbwkMIuhaCXD20+
49Iw1Who4PCdgnQ6hW5SiO1Ns4grZFb0SbWoJTAfRpkgZfN3YRR6txlRZKBDSqyi
Wyq5YtpOt6bCq9rISrXwn+/S9gH4Rm2QXyyVYEhRwwogCF+vUIZOAEKJHW3ECIdz
8xjIpTOxMMuTc7WQHFkWgaR1jbNbnjoVsYK4au2GGRi1Vq2qmoWMwRvl3vKAIBcS
n9zzwGOjDlC9NyBxIiMLD2ETbZHYz8Po7Bb3782JeqSjbQ9DCS1T1CogawdJdM+6
uZ6Un08qKUUkQZduoJTzhrv4yJp3d3GCUenS7aCdpk8TbgoO2Anfeffn5b9u3eI4
LjKNru2wZ9TwhL+FIX+2fFOC/tq6np7xaUGy18c/Chq5JsRTi6mF3XOlhWDmtO5t
YmXSuTExgbsJxrZjYqIK/6vgAtSxvx8M11JDcF7oRATwvxfY4WW5Fqzc/44Xu9HV
7Mip0mjz8orrF3SzETOjUG/jB6MU/AbRVuEXMpxsbk8l8e7C4e4uUOksXI6KefAE
5JffdPWUNF0vpQdAIdMuvQXuvz+xG9KcleT+Tku1g7IEY5nKgqMwUE8rVb5+CRoT
o0vPUikkoMViw4PDnC3mhGBzAXrcmbBuil7YWufBs0s9rdL4zpPKTbFSpjnMzBsA
7dBWhuYsiODL88nuMyEpw1VIGeRa3C5fp4Nlyc5quz0z8ii4cJCnGHdlqKeI12Tu
GSuDdDKQ7C78NSD8Jh4ZyU+t/UB09dqlGwZjALet5r+KnzXypkQZWLKeB2QWwU2Z
88h3I2eMlMqsRhetqU7o/2scar8TYNae4NaAvaHFH5aDqBWKeB4rhLgAKZdNdYqo
7C6rtpzaS8MQVVdeULZ06xLOHZLQ8PSM/Jret+RZHulLu3Xzv1zIP20g5ejp2oj3
UkzsLoxiSCgfVvGrighTAYAkc/3CeSHLoS18DU8qENNMBZ1MA/l79cZWJxQg8qWK
4S8DcwDkGGjbagT4+RNMOq9jcJWxM/N+UGGjwdBa4jKW0qxia6cJvOvKihXQfb5D
3m1oBPk2igG21nwuYkYGxN5YqyB3+5ZvoKxY+fz97q9x/C2ku7u6Sg5gYEgR2Y5+
URHR2iqmmw5QR5Pgc6X6oI8Fl3Yb2zYBtwLUOmgB5OT3MSzpVLLcZ5Zu8B6pf3N+
+53nHewmBK+6YILCb4sN4exZq32XE4b63QH6X6svEu2ZJshYC8Z1c26aDkTAOC8a
bkdU3sdSG4vYFiH2udNV+v57Yy/AExR5kQHTTfjWSAnOGSm20H5yYTxNNNBCnOjt
jBf2x4OgKtC4B3xyKeCljJKSAaMnZo5J1mjL324rRNsd2dyF4OJ57VJEeWWxdKeL
/rZC4YWW0deOOcFW3I/HNdTGqLY+Qsvnu28nV/eK3NX3aqMaclO7x4BJqkGPQvUc
4QlSm7yahpzQ/f9Uq9Aq4KazzTaYdLfROEwBIZcPy6w70OIR15nN/OeTVvOKkZz4
ow8Xf4oKKQM9sk9Tz1o//iPQB7ZLbaQtAQbEcFHoIsqnZk3D0uCS1w3VrBXNL+uU
GbQvdkPx0ZxWwIcz15CE6qYMIuaR7td7/n1ywtJIUL2c1blXhrKaKdD0AmcQ6hDo
65VYAE2jdUEbjYAjauxg5iQ/7Pr6FJ4+yznIeya59srXXBBWTyOiSRU1V7TqZuP6
EIP5vMCU7QJ4UYWaWEw3+ygneEVmVhyd6RsK/GpqoKXExGePN+IAnvwa5BlnTp/t
2bRHTtR9Pbf4aGY6xKZ+RV+X8Wm4itQ7IvRsBvUG81z+1sgrMKdgnEFxzFceC7mK
XVpFmZKcVwA/kvbWJ4T5aq/g07aQ3vEgcwn4aboD9ugyg7/R5D7k1JJX0JPFkOzJ
0eDesKeJ5kBJHvrFVB+FZgtcHS5RQl8XkqybQqzN469UqMSGdV+Cg9Bqd0zcdCsC
ocVDH9B/RLIfE4QGPbTx2bNts9Qm68cmHsdsMN6+pP6/Y0EvkXL7WCOCn5hwFeyV
PvXEGEwpllEwsrWSKcRGvSZfycQsBywl7sfaBjMqNTJn+HzlUzXL9oogKbLkn94v
Y3LInhqfvrcRssFRbW9uycHENbLETuzVob4EzIa9cKKcewIq3yObqzzuKSfYSUXW
vjuNIIDhLVI+8HGKRc6IiBs93JNBwfBkPJflEQd6XSFKQ95eAAOfszKjhOyP2QRQ
RS+O1gV+NRccoWE+tOq9fTT3d5hTtv410WcruJeE0W0YbbU85wN5jvQYZwPUlrwc
TCV20X8nqd7Ny/8/Ct79Cno0Taik/+GC1U6xksfo6iEQQoGhJfxVrvsbx9GVuNvP
qMb9ONKRHtK92ww4quLlJipHub2d8gh7p4csWssMMgMtmbOFFA3zZCWpD62Yg0/n
V+FkSI4I0p1EKREHvkluVSa5pOUOAEWzJVldHjy3rVEuuKeXYsYwB8Jj51kUKytf
RkI7T6kFafVItQJJMEJUhi9WPplZf3RnGXWhx15h0nD8JqfQk4FJTfhonBgXLGaH
Votqa3P9zmsYD/MV/0hdoF8RLfh5dWgdYY4YMfIZLQBIZKJoTqGUusfmdW0YQhlX
QiqiYFCLSiRsWtuyZzCVli6q3D3kl7Sb4B/1/917g+lrA08y3dNDxFUQC5QVi+Sw
7pHfATKVZufiHL7QuXvzjuuF0IlYpCeKG9YsFzZrrr8FGJMh4oOXUdw+f5b4xBPY
fvuxpHI4MLNzoPsUi45jCmq0ysYTFGaUnAjGJHvAntgSYdUmQo1rl2X4har5qpO4
TXdcJqjXGTL/U7gzZGOHTLi1S75zY8gsfoTDUJn79E6Nug7DwytIptl/wIZCuyYP
CKxvY43rbFijlLdAZG6Z7PGo2srpFxKa9TO3A3zq24+NErDPVKAbHwwOfdO+Wkkm
Hmka4icFZcoX5FWL4S1aJfN1v0IVD9Dft3Euu2rUphya2CzymWPI1gSl/OoUKMK0
z+xvwkfI+8Mk/dvpNHcYcLo54H5fVSgdYT3ESf4d5Dwx0iOoILqXdXL8DNkk9NkJ
dN9ztzbGvFpBYUcMObfT+gh3h+jgo7E6vZRacDREqa9lXc/XMmRj6MWuCPNuuumU
lRjrM5pkEydRH0Wbt9PKGiTslB/O9zLxVS1fKpTMgxy7tDX88vP9JRgBRqSN1uXJ
pqSP6sbpp/2x95C5cCgdOQ/TJzH5q6mo9DqFU+2pu7sFVzwV5g+BbksBhb3gs2aM
wdyaQ+5EoEu4hap0j7VMGcqW4pRc75VHCvQ6dK1cmrdqdLvaBAHeLaMfgVOSSvdv
wuTd4sLi11wZxpUBaORxFGe6zSFRQijjyUg505JQGOBnuVSx8Hj9A5lEs+GmtOXU
JIzkNWdWM3JFtWb8rpyRutIEz1tzo6aDm0AVR2dEdEn535dlGEBOQYutMgfmfh2j
DPqqncsPE/kx+QLV+nLE7VXFB6dZU05vuP6l0MnqY8s20jOwVzzPPT1jM2erjIgr
tJhdC4waBMoWkJR/r95Axl2byHVeebbdfGABpcOkpWG6ekrQs+bptKAEtyBJZwjv
FLQ88o9cx73TfJCK2X8lPcZDtEA1z0JS8FRMLAyUQDXKgZipkGDsa1QWKpNPxELv
P7RRGkXRk9UvJ20gmS8+z9FV2JLFpC6PIhsnXTMYr/RDLO7xarnlkIGktgUj1578
cteB6lLgHzQS7KKlGu9KOke6D08HLYI8EPsCu2R7IGBs1z0xpyIROi4WPNbyDmJF
nPpyp4opy+mljz6BFoDCCCTuapjIp1JQL+AUnLBfRyCIYx7qXKAVWUi+nLLc2Lsv
TYH8WArQx/q8YRQkbXl6OmmDN3fxpLTjMqB9Hz7XvIiZoDn9NiazARdrr7+pR+rJ
FPtTkRVmSYnqrGLORujjq9n/sAGEWKXitcx/o4rL/sOLPagNFuVJE+FBterBJF0J
heoeTa5EeujGmog7Vl/Sb28jueje45K9uIGCbXVItCUat4om2CQdHPlUJmgZ5rSg
z7HpKEJ8+o/ldTLjHJQn+V43isZSMwr6uP8i1OQ19ouOYTsrgRvR4po26OTr30BG
MbVX/AnobPsGT8kABkNnvrB6YTo5OxLEYnerHrZhJUlVoO+tcs9ECLRWZM+SnByC
VDeg7HF8QXIifX3olTgtVvKqmTf/Dg8Zf+zqwdTh0PkHyYRN6UGqwYQqgR93aPPQ
oJkybycPwVbffjIA7tu14BpaBlpRnDyNwtuRsE63tTnP8c9cMg/ss+m0OTtYFane
g+sBteBPk3GlpnjbPgm6ASxtlxO5mP0MV/+ReEWaE1WQ4FJ+H5Wksau2QgkED3ao
rJ+PByrkn/OZVczBCtT7NSYq6kzzia9yWARpK38aHPYk4UTN9jIoQTltqJ7zBpw6
BgF1dseEpN4NQq7DLAmPR1vIjFfdOc9u4c0YZl1k9iWiiRiJmh923NOl/KuODsh1
M96J1oMyNoR9RPoHSHqIho+phgLwJ6+gEJDqHkg7sQ7WRr9FYyx98r7+1LuLoOuU
QJh0r2cYdPI9rUt/tpzdP60SBNVFdO5VCiaBdgg1f6jJywtqGYcoYUuQRgTyPWG7
2whcvcroLXeOpe7R3bREzhmv4ZXgPjS/vO0akeZTgZZl5oxqsOv3EC6wlk6wGSBp
peCg9sBmndkhLd4fYoCKlA76Qu5fER0ixy2WZ0v51JA/po5rwMMGYj+75ucLxuMY
Ru1h+ayY+K055nRgXOnMIuWbrPOZgPxvalSo5pysFqJHUB0AF3YaYUbdyqXtQ827
CZ24GdCNZXWmmBi6G9qRnAHnOJ6x00C3sbUJyruRq2ImAVyvuyXVMPdWelieea86
8QcmV2DSbLLaZpnMW9+Ce8PJ9tkGYE9q3CsGyfEeTcCRon6wPpAi+aC/sm22D2h9
PmJsN/4ASAEV17z59/SwEx1e0IYUEvrPjqLeLTwDtvsktjsfWAsuxgK+C42nQlBg
gZtvsrd2VOD+vnB0Upiri9XqKLrd3tb+G24ymNp2+0ikTveh0BT44Wl0lX1mG7C9
OQgmXahJadQOhgPW2OnMD4KBg4aHzyzpNlWPOrnkxMMy0ZlhgGjsUfOiAadrejb+
58mI2xRekO8PE6lkQDmS2UbsZ2nZk/Ass3NwmcTnjNOe0idwkPGtvRtkzbFC8shI
U2jxI16Mtt7I0BRYWOb7okky/ltfqrRVDmjzITKxl3P7M7TBHrNJ4Y8tZvsZEj2Y
3bf2WKuk+yC18blLS6KkGdPwvL4B2taE9X2r+rS4Lm1oIWKr6N9UKNlmdsGfx4GH
QLjN8OGJpeyWuJ4doWcqU+M3tNcctM6w2AIG3vVU/3Vx00F8n74Q5JYx/T4ebl4R
Gz04XK/TUZG3bmcmn+NO4Kw0HP8+2F1jpx7VE5vfLo2i4gBFaa1WrA4b90J9YNT5
c6IscHI9hA/jO37G7r75vwuc5eUT5R42ARuQxZh/gGj/+mFkLuJMG27BF99wFNxY
ebs7iqkBPTZGmrs0o6JCEwDcmK9r1/8n0nt6RFttw2w0s9uP6MQMMVU4b0LPTh+D
B1v2jFrqmnFSMpEjmGjz3+1xveOyPT9F4FddLysbpfyS9NS7s8YIO+08XIvYYl/C
3vQezv8LumuvPh86pNnf6w0HCR9Rr227nsGJMtlex7jL3LukMeKWEn2c9EMJpY1O
XxEnuZ2dPbG7t0XefLt2f/xe+qUhQtpSjLeR73r8RVn3cR6vl+YUUNvnvrsyJ7Rr
MV580aDLBtuPuwgCCyOCHayzLi7T8JVd+qk6j+jMyKmgC7NVqrZh63VjDOZnOGPp
2HEdbVvMbiemnD0UQHp2rvpwo7JxJJKLB2SN6OEJvmHb054Djz9iN7EhjgINIgFZ
xECQAaLZ3ikL//DPeF5iEBYZ8Xv3/1o11yYNTCNc/j8k3vKHrVKxf3wngxbrxcO7
NS6jfzLahEJHsH04wXkaj1o6H+Hr2WLvse1jb97nTKAA8Q3G+mFKpVxnT287n8+x
vubqtd6t6PKAlQZOZovAvmCfTyzIxUPT6mHhEM25sjVGtqVNu3vASLpkvkSK2TxK
sLN3IvltdOB6+ykn3APzaEnMsFBTdpCztUsE3e5enoNfXZ8YsL8KiISzpUk0hU3t
AZ9y3AuZVZ4QN5FopZx5P0OUGwecXMqD2KBvwAuZoKODFm/BkxDlThxc74Wx/KVB
mGl+VSTgyDosU2rfxNZNVHKkgPdeKX89V3sfSyiq0MwYaozxrlxC1WV1Xuh37JBr
vB4j4Hon9smLcNgU6kG2SJdmx5j/5O5sfrWQKbvg9vgGN+QGOJtaDCcN6vaRyrjH
+znvzcI7ZjCHtC9QAN3FQ1tv9AP0hpyQieWh/3AHlxCZcpgbpKd4q1aMSZ5Lyv7X
+C+d7GzflL+GzJiR/75lyhwkW0AA1iaOaK7KRAzdkvz5URbayNSx/0Nd5swHuqFN
jZnAdiUF/LLdv8ParpiMd2gBQ8SrrQpwNkNOBwPTF1J/j8egSqdcxhTIsi5g8lU0
/YCRU/OKe2zG1MmzUF5Tqj3E3GusFzQquYtuvQt/ACXZXe4Gcq0Ko3DjH0fy9n98
aIuUtTK8DjkCu+HCXlQocyNZdpdwuSW1hwESZsz4e21bxWDwn/+fADDsd2KH9m0a
Tiq5MDEJKthLspOzK345GP4mc+AGMXzPxR0OtWwQ5A6EfRibzSh0isdkxo1yw298
v69HMMc4KOtXFXK5i6sG4Etjn3+ql1OW/2BLZXEShbzEv0/+EWnkOcHKMSLalYvT
Xse7AiiAoF798yGRgkAzTaY5SjFUyrdgwloMyJ+0S/TfnyhzdL+CU/XW7++2uuUH
p7MoxEO4jIyRmh8D68fMcfw/z+oZWUl66B22BASIZE7ANvX+tXUD8tvSmU8u1CVU
Iv4ytNzxpbJvT651mFwoLy09uL3Tf8HZSEoCau1mYt5pcI1IRQuHs9JseNVqTfWE
ghmFueC6sS8rK8wELYNaIqlKddzTIXaXMn6Hlihra0co9Ebw3s/1XB7Dd0ULWXkE
+RPYELqRsGEgJphEs5hoS581HprF50w1fs8SB1e1/AC37B5dQ4oNvk6rqJCcerZo
JrgX2SxcYz/v1lL0Fmbzr4fnsXdOtLurbrV4GtL90VtGpWGGd7hq9N3Xs/+/uSvW
vzClu4urFUc2QVvV2yhlzaRPRviypMnKqJ9ZQ656JTzaRxzaXnAw3WP+K5JEdymL
cmgRUy+WziJPlYSfMBtbaFe4J3Lmlb6AwP5G3xbIbdq/9dq6gnXWWgyuue38UpWT
FTAvRGo6Ad45WWQBWJBy++V7EtzaDMdVOMjUjj4irVCftfo0blw+ALimy2nSnYTi
27hx4fWSN6XFpqDZc7FydLwV0DVE/pvP7Hl4ZNuQ4A67M6auSSjiftApi3Rgk/5r
wYv6LwNgRhQsV8liDSbGS23BxzlGoLRmD+QRobAwORF4G+8m3C/mAt1CIpCBShNy
sr9pRSrFbXs/HQmgJxAe0cFrQ3zTAM1nH1jaxaAqJv+1cn9Ulxgw4eCMeDAtkNNd
0XXkxX4S13kGYvoVuqK0M9r2PmgpEkxwJ/VJ7mvk/gtRJnbv/+28xZ7LjP27ymJz
xvl9WXkybMGEuAX3bWTgrl7zcQPshH6cUcqiVv6iMl0+dx6/VC18BIEq2a/wNZok
CSXhFJFPTxLMstcHbKTe8IGTWmmKBNpUzijyMHNN828Q+ctvwdtzohYLmHVTS3UU
PTPaRG5UVHrwrL4VCMh5UaRbOMpK/BhYIDdh1fsdt62fAnAA3uwPvrP1MbZaeRZV
ceRNO1gPdMJc9GxLNgsSLiZ5DIFFpWFG1U0tFCEBxJ7lrIwOAwVumklvG5/aDquq
QT1d+75AmvTvnNQyCr+/kag/D2J8o9XrMQjqrZNZE8WwtEnnqjCkdiy2prTIo+vx
dbd7MIYLcxFzzgmJunb7kNtmBYeeiCWc2TMZ6LtdU0DDxf4x9LZD/sdnY5frf8Mo
Ff+9+WuHxW/4qYpuAaOv2i0nsUhLGcHOIexNN6fFRydtsWNmbK0lUQvoD4Hyv1jf
PxjFez3r5I1/tSWXI6FrXuRaod3VNinDxFq1h6ixhGCIDpiS4yZ1mj7Lh76MbcjN
phuNRWAwjueUMYXXvC+MXWheXGzTZRU0XVB078vLrMkiiUbVompv1S6qG0jRKJ4g
16vIUfV2KD41k0MWKgM66akRgy8wlOrS0eVzUcg91KbTJ8EUznN+VuNv0yP8uo1O
iLAXowxcaVCTuPEpT6E7xXjwj2N7oGYGU4J8m7Wl7HdpXE1uEp1I2/yIOFc8cre+
mqkrxtqe5g3t9cP4hVW9axiT3dV4BvHmzcWbNeYLr43YeR4GVcEV7VRNU59W4yXq
cV3NrUQFnVuDIXOzeZ+/6EdK1wdRDF653mJqdnNpjBnRfXhYW4EzJHnsp/zKnn+b
jH3iNJy842OxDuj1MSmqqXfj5gu3gedlZ8xmbXdkETd2T33kljR9Jc4q9oKKwrGR
Ej2U4u2Vm3uOWvLyqxCF02l0RZqvkADZiDZXCER3rbm2+D8KWhxVIHNoPEy0KCGV
xXD5Ua3QKtZXKpgPxNwN+S71iNkDPowKDS9I0Xp0etAXelWMywe6vdCIfHLDrGnc
yJ9mrmULyyyTZfr2IL/CqxTXdYi3lwrQUREaQjZVON4EHtIqFx2T/xv2ZT4a1aBR
1Dfjppyt3v83jUJEYJ1Hu35pZloOVedfob92QGeULM0Zy65ztdKZQ/IY4GK3Ohmy
ly/JWRTgGpd64KfTz8o9wuwFpK+APPzzhr5Gew9MAfVBjc8U7ilQPkbPlBGh0J7J
AvXzAZUjrSPf3xOXc6pSZl49+xNouBR+zqGzvBNTP3D/fFgKBrUvMIEAUA1W9gRe
j03ANjsFqE3u0afhFhD/lE18KaEiFbQAon4Lo1P7YrxvdOQbbYdKSB0LLIbZyFG5
bWdNrYIVvGfpnOvq2iMPvTzSAq0dxE6kA539p5DxeKZRpt9nYIcguTBZglszVT/J
KA4M8S9GympVA4YlvvqaCf9wfMU5uR4SJ19VGlddAYXYIF8VMDui+X3PCICMqmp7
N8YGJlYcsWhNOVkNo8Q/SEXMpkc3ZojxGbUG+86ilfhovaOVsU111riKd30tr8Uu
n+k3FSw27BbHpz+1NubhBJxB1GmLjcr1dB3EcyPJwgy2lpLDdjT0aNy2y/uzPY/b
GWC0Vf5DiVI/mqxxJvwGtsWHsWfRziFcXNoufPfNbCa4sfU9ULmr1/fL7qAT0KAt
TZpUUNUai9yonQkjRey/DOKbkWOVYl8yIrzIDsdz+Y9cawcrUsuMsQzDif/E2Dvy
4nOwLn8WFYByUxqNjSObbc+FCPwnchJ/yK1Rv4NeUwz/w02ffeCJgUS5NFNdw0b1
zozNzv19BV2HjMou4UqDCeV4QwjCmJKoTBWvzcef4qfC4p/i9Q1870dP/U0aSjdO
xcosI/YqWcWBFy6LSLvqhtex8snRK2JE/8QRz8MfQItpUELf8J6RXaRdqm9ylXBn
uPd9Of+pYD3rIDXccLvaUkeUdlsEtlNGnu3y04cx+NVurnBulYOhAU9MwZhn44K+
ZRTybclTDrhYBGzHHndWOVXaTdMqM1MnKgFgGiBmOiKztABDM/Mu15CzbzuZMzjC
0PfmV1LqNZYpwDlBMNzb70wRK6EdpTz19PSMQ9yMnGTzXL+r6aq5YdlRQ06rhpN7
4NqcIYcjdwMTi8CCOcjaWosbzUNkJyd/4+M4eo/tT+WkZABBXTvlLtkk4CpNbBkD
KAhF8YIlb8gjzBuME6t6G37syJIE1VGdveHo5TtXtx6xfB6cVHiNNzPWys02uZhP
qjptipgzA/04AGe1N4llN8z7sDwqbOVCMKWYGCmxJmJNQJaED2veyDcdJw6Sui8J
Sqc6UlIoVMHPkSjxZaUWWU6IMEOVr6w6R/Qr+IGYu+esxW9dqq9XFOUe1zzh8sqa
RZLcn9RKbNlWe9tDIOcu7QyfkS3EjPhkArbgGgub2+AdGjdig3V641OF5GtlBRUB
fFApJps4fYYDhjj9How096BjwwYGuT5nqQA/hptbDk6+B8TdP7xagElO9atpb7rH
ZeW0pSqbNu5ivLZGr9d7vCM9zLPGE7wJN/Xli3r3UiDZ5pnhuBddPn97DJg4C9y0
AkIn7zcjVk6hHNEM6peXirQXQHCXRvDWLw4T1kmwI+RDAFkALmwzeejalgMYIelk
EAXARSYrWBn2yyIXN7G0+25F2s5pRQct/v/JvYvdp0diznreSSrBb+hOk/CNj4Om
d3rv6GC8vtpd0ujDqI2ZbT8nxqifC8meapBl8wzR92LQLT1Q9Cxh9Px68kjXEhCy
+1q6OVFXYbWsLAWTC2balhYTE3Xjx9JLALANu2mpGLlfz49sShfZWH6U/YyerD7D
gK4AovdRx3moI3J/VcvigcUHUzTnJsp1KHcLkgKsT09JzhPXYsmd49WcMD+xEqUZ
2EHAUkqSPXoutFXKWgJOqHb8SjZ0viV7X0EWiOrf4s5du7lpUL8bRhH7QRa4/crJ
Y45rqHTWLkct1QdVxlheMefbyc9M9ue9DQx0cWxKa7Q+fn0OqHFdiMv0p0Rc2QuR
tc2Ig+d8CbWwjLexktI6USollVTgRQUvoxKcnYBZGsmq84wY+IypDUE96IdpoOxV
vylHBs6ADMlpQvwaNLXIiq0274aY/RA/03NKurIfQLQw+W9u1O38L6EH/eTrVB9Y
I9aepNMDOy9dF0dlnjGUAgW+hHRfT49JYWtVvCS4r4/Eq5UJ8D7d0Sal9wuO4nQt
fWYM1s3fSF+4fR2jDFtycp2N7pi+GZStcEp116HcHGWZYtG/EGDxUxOeNH5YGVNZ
YjxITraR71E9Xk0OJyHV+fbb+/ofOGb+7dlbExSznLiTV1xKucd+iyVq+WlFvk1A
lNEY7Saf1h219oJSo+eW5FqjR5HFY/ddYZpDnsxasidJ++dMaV0qPOY4hV1WGY5k
C21Uj5jHxjgZgCfmdo0FlRdbmnA6msie5nnBMz9GfJXwvQw6z+jMaznmOj/doKMG
PXGsCZow+S6h0DzWFsjA8sFTZP78xPr/wX19+VEJZ4PfrtdinFIsagh2ljJPqoBW
ZsAm7wyCBCEbTRz6JqBomyekTvXr6+2JAFyUnFBPLFH9O/m4jVuL44NUC/qbrW0o
zJJmCfTRadIrW34lDkwhdmmW0L62RmBzsNbsAAg8UdcYgzH42AbEBxO2V+0P9dPR
D86D4mmdBMTJ6uu7LKZswZUdWCzv/qCT3NIrP65LROKcpEcQjR0U9FDODf8wedF0
oV+dlqAiQoft6OqzlU/uoNSeJGyKHecao16diUrhusZ383F+nC1qPuWfMs4Do84K
caTq3EJTB/stOOFFOaw1mwDy22i0JhcK1dZAQs7Xq7/WtsiORZJZDM+wf+4Ck4f8
smjop8O2Bzu+EhWsMOawNy9VKo830RnTe85/k9t8g6d0LUri3OI4BXoUDtUmmkJg
ndFJOGA1tPCgo4/7TAO4CxSGFUwDBQJ9d295eOh5eE+5bgV4iOWYsloVOuWIa1sC
lsYARurPC5a/5IPjkDVHR2m5t095mwUpwzJeGIuI3Mdjr9/wY2TQgEyREPOV+/AD
PF/5G1XE6BUCCXvBdgBDtEu5Z8lUy/uQmTyZlrFHy+bR/hjV6HDCe2HQJZhrHli4
8yUt7k0JoHYC97jNmLmjIOgSN/hvYd0jY0E93HBuj3+9EtwFr+T0MV0DfLzssnYn
UK7VHIOPxRrZ/qVUSDT2ZKw3sk/fkBqIxbxlfyVGhBPTQ0IferLuaycq3GmIh4Vj
I8qX9qrz1j3djQumLrh21OOnCGtE8sXcj1AIhEHviJu2y5FoCBPQeZA1G77DSYxb
LqTGRskROvyii/TxYCSWixX0/WwmwSBh+FK9GrZKnBjhIOQzxBWzq6IjZX/2prXt
13mX4HIjJuQN76hu1UVToYGK5f2rjtIN93tVlphUJMwnn9LpDzroYtq8talCApfs
OodRuL/xeACIw5fGwI1/5798zVXlAoDjo2jDDmgftgyi5qVl5U5qUrLP0Sni5Hpo
hi/mRAXv7l+OJcHMa9C6USnw4pSBmm9Y846/G8eMhx7JDYXFgdmj29uJ0bbi8LV+
v48o4FirCp2O0hKlcf2kn4Ll+24il06BiXPmSNGpqdF2FcljxhLmJmYZSgcJirKy
ttXJgZtAu2B4gRPZzC/n0tmdTGAfxgoeeyCAfvBFpoJRehYrc5utL3Y6/ZWN5aiW
xVxcAXxKV9HSdzBVcnJO9OzeVNwaCPrgBUmEg+I+nni3V03uiqmSGTO7BbXBBB06
eIEYvI2vyPG9UJhYBEtrFLkcGIz9uyc0BBuXWvOUo0RpGL2/oMuKLr0mzvgwh+I9
A8/1D75XIIUBLqwT/9XpcOG9axvD3P91hQ3LvRYWYold7u5GdCDOUanVS+t0yuGo
bSh4cfPD9ihRAzfsIpuygbY/uKPe9flxUtLr/g8x8G1H+x2rv2fht1dT51toNDHz
whh0BKfVWjNX5Nb7N+aqeNSaqkZrTXeYn/UXFXtoE5hRZVBZoU0Ul6xn7wq292yE
OncciKSbjxw8su5z/m6LPInfUCuWsHTR3FRyqbUe9sRRlC86S+7dde2IBYJkStSH
DmqVbcmcuVEqWDePw9YRw+rPksjsgLQdsOsQGGNbmcoGoMCM3BU+dDqcOjPCFtGi
GeCp3szjA9j9Wd9SWclRVJRv4QhKfY1jnnVOTiS6FoijVUrEUyiCPGOaX4NGJ9Y1
xxfHD8Is4XQxwc/dsPG/Pc2t3BjGjPMnh6Y7zWTPYjkiOQbwKxCdH568DYYWsdSU
BFDNaUsdqVk3/vI/w0c11pkt0618yctGR6nkud8Nd0tVeP5U16uIezj3h6VxAwJA
5t33TU1RP0xrT+7MG/wZ5zY61wBGEPOOq4sTQoiaEE7S2+sKY9AlxzaKasSnf1YR
oXRuAniW16BjUjBrlthhg42/KAygyMnAuLiWuWtUZJow/oNUs/54CVJTgbJ28GRO
iU38UudcYQPgWmrDVTcGoOGCJjBQJ7m/+DBZyCJ28DICtrikYJ7b0bhJpYqq/vMA
i9PcEmxm44tMqco9p/0XtjloxD5joicKys2y2sTczQiKoR6rpyON3vLCwBqQEmcW
9LLWBldKKpkJQcrspNAC1WFZ+l1lXaT/vV/qrLO7gBYp+cCNT8OVjbSiNUcp4iQ7
65IrJ7jf+Kls56v5Y5q+L+/Ys904OrNBU9wKfxv6F6qOssIMTCfvKpPSk3jOOUc6
aNQmxInAai0P4+2aCD4FnvmHIZAtFlUuA89QVX8n+PoJNLCiNouhxxX5dG3Z8FlW
jc+Wv08gaXpJUvhbTeUyy8LOwVaHQLwnhixL0cVb8PbkQS9SJqujYys/QnCYmbHJ
ZVPGSeoyrmVzVr1ZUwjRQK1d510QOIyMhyTXp9Id+rAIs9X6iqOVkSjOm0Bz8KBl
phPoqH+xPAXXFVQDxbyOToe0HirQeac58+KFKjXCpcIxUv8Q2vDc6ZZ8NKAmyYFS
Q715YJ4nhvoCMMnIRuzTJXPvWvbsuIJIMvFahcXJC6ewi6W09UCRwbDHE4hP7fF8
mGPRkazlu+au1SO8oRPjxoyQ6a1Wf9j8iuTiH5K9G9s03tBYXP5FA7ahdWVlt3HS
ZAniKhWBNtykxpT0HYg+l4WUnJeA6fDPJKCnnY31KW53V/ZUFU9suVY/i2he0g5l
ln1THIdOFUtz2lLvFN0YWJyi1gBxOGI2ozP0WY0G+pbZMXNrgSezbvKkeXcKNcJT
yVG8UqtISac7SnVNw3e1xbUoDRdcmTyPLGmw927gZ+6DSrE2/Yb8VjCjmTjBcuiz
z44hMhX+EQZBJilDSGCSTZUklLuZVpdOF1soIRTPSvHHELFarJ/r865OXzXYo0YR
L71QEwhG3j2Wmp02SjPIiIkngyIFRYMJ39XjOGMGNGduzgusKurUBiMe1N1lWMUL
c3ugAWNA8+IFMUryqqZj+5jMsH4RSmkfUPjbtJboKfninTK9nppClf6K58zsiEtH
GwkfGAeyzt4N20x/2j8sjBl2NWk6sbc6UKZP1Gzl6sHY1bzAqM3hGSDa3uGPMXqa
7cUqc4Jy6MBw7YSqgKnlHM4cTrQS+81Pp9Erhc1SCXLOyaG5q4pHEmGe8QEpeV6N
CfVXRV/285dIizpd9xcakHP4yHWFb1eBNeexucrFq/cY2LTTfLjP7U0yBHDC96d9
Os9XkTJjCyldbpJwWINF+XeSxFvlrsFl1u6Reo/F0rHkFVAudo5fV7Uokx4sqeZx
+gNTpDrI/qycEtOTZWLVyOaFN3aIlUGUBcPp4BG5u12ec9OykyZZJqWdJatjMTbo
MM1Vj6UYLHo9TfI09ZctMN2Yf6XZjOIbqhY43snpA8B/to7mWeGSY7H8TOhE8x1V
fZwjYCb1kkcxt+zW9WAmDpjgBeEHZ/itwWfbho/jKRiIK0GeFdUynW67aO/BSJs5
qR0UfY9yb8qG2YS85SV+l75PqlzD7vVynXk2ddB+OEXJZZ1qoIJe7o8W30cx0A1h
RQE/wLEt+Sgcgs6PgkXOP9dnJjhrjhqqhj7Ub64AvQNMnkUHUwpbeFq79e8OmlFp
bmIcaW4rI9JN0gWAGB4elz+WPX3PwtEvSay+4Hx0XU50JTM6R5jibm3K0qoQ4h8l
8Uc7JwZMtdzSV9MYNLiInSkpgfYhguMBwFvDy/+vV/sDZIgxG0tY9ziIh7QNETV5
j9JDX3c/hTpian03hDSKDqV83dl+KsPPGMaBKYB1Qf4rIAGu966urh2lB5Zd/2/m
9xqOGZeHzlcsUjz3JeQ11fXtZKZAgHyhkEFkbz02weZlwr8w4zT33I8D9FiTUY7c
hDMs/e/qOPPi5YDGrwctCaK1bosQVfAqKj/tqcLWVqLkYiPGj3G7gB/hr6eAWsqU
IW/pX8NOdsYbA8cWquCMRU7VjJPTCfgRMEnwJ9su0+qqYSpE78QJVizvVhUBBNJT
shlA+BcfqmHX7OlaBPh2TjHBuBPiQHlpxDrIly6rpI8X/xpTgeEeWVIauiZLJmZm
8UTm1EFZISjHKd1OWT21A/xHA6qoRhxTVuMrsiQjZ19dwjzKLWVmFYj2iImKVwPC
idQt40PZCe64Nasamy1kAqPenoRssbXDXuCdaDkw8tYjKUpNqgO7CzZmTIeBMGEo
d+4Jj91w0RlzVabDJiTN6QfmVCiLx+S6R/atLdspwd8SW5JH1Q3PKK1gwiB7ReCW
ZjVZq8lblM2cjVMx9PERmEzJT2kEAw56y0KRbQ8RCgxgpYP3YIfOhM8BN3J9olx0
52XN/u+qjV/AezcKneXks4pZYor/7E6L1W37RZwxKpeQzoQEAJtu8eSLIpg9u6xX
CJN7RtZfnpuWIPP1Xz0MQX0bbkQcva3heliU0IgJ3eTPaxSSytJARtCr1PIFXdjz
OZj8djtoxfSCPfv0Sjcb2ewlg4vgtD5uhXKvws3KAPvDqyTsrGXqAqvmf5sVDQGM
shoBrYaUP5ZHEKpzRWrkaU/NGDn3fOtsd/Z1RNhhNv4J93ZBy5HmDhWwMchJ2mk4
otl4qhqUbOmgL8eQ6GtTLFUFkCxVmzAa62pF0hVH8OdED3RB5sPdQHCMg4061+AZ
M7jFsiN41jW2MOf6ZR/GV9sTUHNqQkfKKABteEPVDnFLO23Rd3jUSoh/jLnAKrec
vEplWs4s6gIQxwVwm1pwYV0XOTSEdQJz++I0l5vgvHrRrufubJjO6/mHxQu+8ZUG
J7E1s3ijTpsItXFY/kcxbH47kGPcw1meEe5Fdvo34oGiUB+x0nZS9Fqqly0Mw86d
oqAoCVUY1rPEAVR2Wn3lF1H3Zq68zysBGQ5+r7/d5g/W5zsenPtYdUCWwdM2UP24
wJ46AV+q/yOungc3b3r1JySxj2ENM+iaANNyrCGrLzHnT3IrsAJrygZQ5JjXl31S
02yOyC66dPYphl0AIexLmnw7aPF4r5cTzCcY4cdZ9QYk/x+KeQ/nT9nwGIT2Fkgn
FAXje/RcXlN3AHfnEzto7byhwAOzoppP9GgGilve5aAOs3W0zp05smuTElKvHNe1
RXopGY6tJjA8/Brq/VNKJtUww/9bhlgo0JOYqTI1NllbOF2IZCYoaKj1/7nLe06u
LcKQZVGHNCdGTPrUrYJYuiBGcoGyJ2Vl16davmdA309iaF8u8kG0UB/LOW0dXmA5
IVXDkd9AEwjhQxIEAmTW/RRw7/jBdyvTb3bgLJ8rMZyJCVmuSSFJKN+LWnbIbvOw
1ExbSeVEp9m1oPwLwhWxQN9DsU3dpy/AblCmHZBFG7H9emENizkbtdpvX+EATlGm
AefF98r0UV45H2e7p7Qhvd10gH7yxlfLWH1uyTbsd7S9delOL+nQX3IbkLEEm+FX
jgTE4+RO+yts6OW0TrKfDmNBwK981/Dv9L9k+oLwjT8Q1jgNEt0AKrRw+aw4NVH9
8o4npAtOXtUFGd+3OdEjTa8MDIzuyfoBcc+AQsDDN4+5TZn+UfLanmQe+ZM6Yy5Q
z5HNUCsh2ioepuqOrtbDAr2y9iN3Pn0FezOFKby8MP2Ch3sF7uDI6EZna4nYwmdA
I7wTeOnNmoMYTM+oSINg9+eG39AGIDeqsMRBFPcJzfWlm5/q8mXlOmgZMdYeNOyg
8ZZaG/6f5bkax5+7kxr2JHDXf7lC6sK71lnSuE/g+dGn34kiEY+6VJfkrMOiuktX
xfiZXnZvzxs/gp/4eosg6scr9KyEMg5mS+v/83Zo6MFT6BeN+KgQD5G0Mz8a6au+
YymyRd0OU0f3zyHr8EoXCRWHR2BLwJm0JwY/kbgziCIYKi8WyZkJgq+gZMmmJ3XQ
qtrn6dXyR/L4PdoacygZUDFP6028RJoADJ320OMGvk2JMRsRG7LFFRVuaM3Od4oh
8tOBo+JsZXBZRhx7zZsN/RG8dbvs8dUVQRr0WmTb5KSw7Zxp2nrti0RaQt5ZHGBV
A1FQ97t2DWWW9A7EEzvtlijikK6aBrceecsDQo89/IT6nBvNfXAtp+qays1H8qYf
3inMPB53T1LYqNcnSs7OjUldDuz1n9ibhpS46aoxGDQvKDb0KLxFOgvX5dpE38OC
6kUfKM8C9diHQC/Hm1XvLfXp7vIrCjnr+tnvEoA8TtB7qdUOlIPQNeF9H5h3c4sz
8SIwHTu1EXzCmOm/QGskGlRQMFF6MHOeMHSKVseEvD1Yft9kjOC/gL2Z1lrBuYbj
RehmJwMO1QIt7mEweNDHB+hsTZxca2d+5/Zq3l+ku/BxqMAVRVdy+1PK6TR8YTDk
i2o+dgFWZjzB3SHLqDELjbszarMa6y/IkU5zZeI4Q1Z3Wz3cq/L+FXdNClKO/9ki
Uza5m+H/lCd3WWuyN172jBw+ZM5iUPUxnBzWilxEi6cyiLYhDz1ZRkKnWnleDPj2
9Uov6IPekXakdMrSsUDLVedRaQvw6dZ+75Oj5GNVtKk7c9Ary9J3ezV9mEdkd6QO
7l1C/AwSaO3MyV1AKCHUk9AMyI8VS/DZ6yK+sxDWqsvSQi+p7lKRwHx8iCy5o8r5
dkRmFhSOR/PxOMZcQvIHq5Mz3LNbeVRgzC3872TIkVSt//sgJGRFy+ePf0dwZVjU
WvI8C5XPcDavrlDLIajUqItoxfCU1gkQjlkJtCej6rjUfC2apv3gDZ8+4JLHkur8
K+O9y6kb97PhK6QBiXSApkglBKi1fNcimJ5xrLVpZj9cW+PzI7NM0S1ZHBwiks52
kcYbgScUdWkpo6RlqEgoCKC6syVz0kF4G/Y7dK0MQsfvLiWfX2ePe4pqVaDPYonv
aTzxKWgRlODdxNHK/9isSoCak4DmjpxOzpmJv2zINDEAXfi8PiEEcUgj/4cJo1Jd
+T4PzlQk9VYqKNvrsDIYoQPaYskPVhlx98wufn+5SOTYB/5l3va2Hlzu5Ee88Zmb
yzY/UApHlaq2WPcHk1HXNKVbdRSzlzxCy5gl/WZFaGsphfaMn+h5GJL2LQ4yyslI
sl0UmrM0vnWgjP+ClYDrycU0auaWVfxG7lGkjHjVJtxfHOcxQSCJmexmInufGN01
rTXpf1Bzt3UW9/PVJx7R0tgxdOwxasZWQ51DgMZ3SNuSHFUXrx9dIB2VeaLuNZbr
IHBsRdx6/0WlOlgok30RY5abyRJvRCBwF6FHYHXEzjBT0GsUP+QK8Gv2LwTdXsht
Iyt1+b1JZA1Mq7+U3OmyfAbHtyge58GJeoG4sLI4YoBZrDeBHZNH3Dgyz9YWKQ0E
wmTCZzYNVXrrd9lmy8G1bTXO6l6/vUq66+FIRs5ASSMOo5DkQNEG3bZR/7Y194qZ
gxWIEP+/0oVdPXSyFsVWS+AKYbtEhPVUSQzussBvZgi9xoBLN6781Zg66FRPlc6R
TGfsV2VdMiWiSZ9wM/vViufSD8LV3+ndzwSa2dWoNq/4THU9758LEg2KZr98FjyO
Zxrva5AZN9aJeE7yNP7VakQetTprDeFSz9Y1os07n5iDhMU19aNTKbmXcchFCs6+
VjSSLepyDt9d7GLbFN6a3oLaPN3ApAH7if8rBfAhVB9C5FQAejm8ATnC3JmZX0oj
8N5uepA8FoJrWVJAeyS01z5e4Fs+dsK163NEy9ZfpFn6Kl5czdyT2SNrYn0iYMlg
oz+G9PSXTzuWAayrrj1Z/boFn7RNScpdWKC2hXB8uIcR3moz+Xv/S0GKXLxCxOkI
41XlTaOwZ7mso6jDbxzd851Gu06MSC8+HLsH8aTcV+HlvTtGJd+tcb9tdu2PNFKb
nNwU7woPM2Y95DhLLFPMxJrTB8faiLQII+g6drp1Dmc75Rk89G0fYeNk46wsUCaB
URW3+XfnVY/M+fUbPQzv/Te2rqbRWgJiJ3Sz0Qyhz9oVoYwSuBCChJt7XwpBnSYs
CbKv81yzRp9x/smIeC3go8ZBWD87cYj/6Iiy7+2t4llVL5JE4IsYw8b0GAZK9hU5
sH3mstl26YudhAtk+1QQlGRcALwx0hudJfHEea1y79pxzt9FEtxYKR3NWcX9lr0k
MjDb0eeV6Xf8VyxonA8rfDIp13fTfeo1WMA1OfHOC0GEGep0QNbCsnZW9LOXRPis
gjR62eniijWRVjzq89uod3B4Y8LatzRA11uYofr/ulxKr/CLlWgEzcmAZW7z1fns
VkDPLfiY36gItucV6i2hCJOgIQvG9DQh5CZ5Rg/RHfRMuRPJuA2bMl6leEcBFGdo
q5dljQhzxYsb9u+JmlH0X6Woda069lE2NYq9AoXclP85vdI3zj8PUZ+aM/dwBPI5
0M153Id4MvylNdMOGfH2Ep44xttkM6mk5l69kDAeWs0V8lVxMwKkrIod7QdQehmR
baFEHExhbTveNFCEU3Eyeem+BFDq6qBtksijOHq9BnjvVU1unxyz1aZqVZ13Yo9b
giroGyAgA4ClBmhSGUv5FIydmcynLJ2gpHrTrzGdbyIMPP5Rujb/q5EmjBYm+XHO
suTdicdC9q1sHcXEhJaBxqccovL5XME/0+yQVUsKiWOGDz+/96LMcqm06rs8rnym
+SOaJMYXEgP+kAfOEjy4Py2qPXPQ3/VxCRCjmRn5NgAl2s3Vou6ENcJnuXHCRqP0
ZKW4BgBUqzhfmLvum+rY4vpahZae65Jt/FbcmX3V6JWsXkHEBmoTbtTAAH3A2xzg
yNpxI6yOK4VaajHHfMzJ9XjkRN7Z/z7jaRWaDtSNPELSqUbMPi7opbZo9zrmYG+u
b/0tir97+EFdRh6HNbBd/s7lnpGmrBMqwjHYxSqcu45lmxyMnVJecoy2AbqQ3OGD
95f/u1s/TK1WL5anAt8Rv/F0rAN0aPUhWSyn/0T8OnU2xZhB3pVgPGtPTCQIr+ql
5+AT4R1xsNvcRx8z0LFlbu9IpLNK8IjI527jsZKUUb7b2Ac5Whl/KgPNRA9Pm7T+
qDXuNXw/LaHh5yGZ7mW6auAt8UIq5SqT9GvwvydOSJPRepxXgAyXZ7uRpvDFEzhf
N7KnvIv3FynCg548X4mEOKOv4FcVUWOkq0YvYd+MbDwDGf1rZ2zpnMQNLUgUqG8e
+WZZgND7akysQ4jkDGC5JfO7YhamUzDnohcXS6tcAo6HVj1BPUVFSJ9kjOPpW0i6
niIvu9moZE5MsIelph5ycz/xU/qgI3H5jMeZg3EZguXB2imtqhcrYuyHVzk4DQjH
OM1IwXyIEGuP444zopDa04WwC+Yr/LIfqMMERZ8TvOcdUdxkIiuWOsJTtwmYuKxY
N+8IWPsOPT2JjD1OOaCbnbYy24f1vQanmK4whFNP+/I2e9m0MXEkQV2yInEMCZfv
TD07KJP7JCWu1Sxm8uu/VuNbvoS63VkDjoYWtoCs7NeQkrhv23qrG8DSwjagPoXB
y9z9yT3lwKFRtmGg6D50Mvo28y/8GLDEBgFkaqCllcLEr044RDhYg0iRW/bMpZVV
vS63mwj2LQDTzvGYadZi6scvo9zxpuAq0bOSZrbfwEssot1BI5fn3w7dTiWGKHIi
g4oWtOcrco4EhkZXmwRczY16JGxVzcVeCPOfWOUtK9t1x9ZR+mvHwrLwRARBeHcG
a1UzzMHZ4iQhLg6pJjIh+goNZV/5u7gMDOxx+JpVFf5yRusp63D0ODClAKKFUsVA
nHuoVQJkJuMByxdU2ZV4y6SBXQoyUeoT3wWgE2qJxMlPKd16vLwO3i2T+ZRRU6wZ
BQpiqaCAvtKfbX6Wvr+/j8I48knsHq829JwZss/D/QZq2fJI5RKWY4UYrQQzniHv
XLtjfCi3pZ47y7NQXuH/JbspehoP240XPg+F+F0oNKG5bj4i0ILHmvBbqeXkrH2V
bbXbu8k9EBgQbDAkrxrHvX8c8aYuwIMrVbdEaGFy8IZr/umkQUVwlmublAxGxa7E
YRrfP6gs29ERzNayXv09tPipmspG9yU+fyM/oN9XL8S1AvqdaD9J7qupd5UAqphD
FUsvaPR7wn4AwqbitBxvQJS6IYabNNsbcmKkVapzpZtuhxi3AzbbGXvQ9bit3UXW
IX2YrkL7G/8f2KOlyan2HcLrN1Xhzw3xyfY3XkaE7EbltBCNIVjc2aveOabBRUkD
1WRJXyUJnw37uLvOCbESm1xVvcwTU6FxePmLCY5dVNYA8WNR9bKGMS9BrDDN6Phg
1RTqqsXIbRwYx/86KxEpZBHK3ocVWI/A/1KW1vaJCzRA7mmyXQzh60jAsVbS0Wzq
OPUKzIs0hKo7z0ufEMGF9LhIL/77gHE0I088ZtDeaf1OS6QK8+PrArLk7E7GxOot
wS/DiZPoPPrXhU1gwt4FC7kSTahKwP1NXpDsfZDgzQX+UZtoJ1WiuuIOiZUm26fA
ifTgo3VejvnVJtISf0m4la9NesNheev+BjmEvAWC53Xdiaydt+tseg13/pdhTUJM
BPAkmBPpeurzBSlTZTaTY5dip0e1Bjsg5a8gkCt+TOUr1Tw0pU9lfM7sbePB+ONf
mdwe7zvWhh/bvIyihSfbpOJpdlRrO+mhAHJED7VLVt4xCq7NclHXYHmf/vyK+dTO
Y9CWjcu7JH7zq6bXw4+ov4o/ky8EXeQBqJKwxX6FlGNquFir9b3ES2eKWaHQ6IQX
hNBzEnJLgQ9GEoCFmNIeKHnNUW1+DpmeAk7dUk0grVTjppjNwVxGzS6xPZn8LO9g
PDoRW03YFDv5V872kAnZxkSCdiywYNgoOTpCTf7a2XWWJf3sqw7rgxufo6/EEreo
t9FbwSulJfCWEPm28zxCa7Czr4lcqfPY93IjeVrPvTtSOxl5ZejJIOsBFS8/1j3m
43HEBAvOl8Z1/HzLCz92W9dqUUvo2VkXz5Hr8AUIZMma08iCATNGnS3muT4j2ieY
4lS7H5/323ET1vZ1TrQJ6yh+2ndnV7BO9GY808wTl6FyVllWzrMdz1EJSn9LwIaR
n+P0Z68VbMAyskUxsM7e4opDFAwA2lLyyzlEq0hgCwns+kw2NzritUF0WzJkIx0J
+ZG7cuwetgw4FYBWcVkbd3m+zW0VDuf5HVXdrqmDSqZsFS88aduMwzELCaeMBfYn
KyaeEdGOSbtOryW5APbe+8CgymlbbkYcYLrPhzHaHEOc08Y9fQAUesNkQa7NsHJ0
hKTizDbDSTGZvr/gX/I6f2ZNx3qPnMciR6iistin2XQXZ5lrux1oaf+v/c/nY3Jr
1wndFOj4GFnNDqtKrhDZ/KEDO9JexDVWyIBz1lW+g6v76EV4J/m0DXIBc/DRKePO
YDGlzbscpyr31GSICu6B/u+BMuFg35e+5/7qeISesbS3x5BfbL8UadaliMh7RARh
oP++NZ5cTqWhj2pdP1sjg3/h2dboJmxf6Ve4/fpUhwC8dx6nvJzx4aIXoxNTVAA3
t5ei0CQ5mHmcQHlqrFnaGDXqP+gdvyguM3CLJdwbsHN2PKF/H/+HsK8JJKZu/5Rx
WoqHk1mgMgjKx5XrsDH0qdUlg0Aek1SPCNvW7UmXRi56+54Z9KVaLrxyFWf8Cwzd
YZFQ5RTrQqwO5w9caJugOa/0eAjkU2gg0+H/B0SXpPjqA3JlbL2vuW54C1AkIrrX
N25tnzmnw26bFxUUNb//G1TqjjrD8DJEq91HPHzgwfax8fOY8hoQamstW5gjQBxH
DIwkopufeeJPmIBvRa+BG8OtDgaSSvAGK+gfTDKSpmv0lNW3OILTJVh1mnZWblKl
c/CCVJRJxvVXDDFQN1qeO7lu/l/A/zRJEtsU0FYu2qNoDey+03lpe4l7FR1/RLhm
q+9QP82IwFDrlmELxq9kvM+bHpHCCUTTYs2JkbRV6yZ11PiEXAitoeBLym/UpZmJ
Oa0dG778Ouh2k7RDyoOtH2hgJ0x0euL8VtbqDdncwYVHQjfdEHWJNU9g2OM2bro4
Xe7SJEBJ5gfo89HlexivQENtIw8mM4OM/1ioVEEqu7PuZfQbQJYiNZZWdA2y9p5H
USitJX15/BIE7NH+BWbfLXsZGrcMli11aNhdB+5ccZLXvZ6lk58C/Eiv4gkNZaD4
MObvkZm0Il1WYVO0FuKi1tPTUG6Dz/thwQ5XwDw7mGAj/OLppeK8EQHXQDTzWtUO
a6L1WQKigxa83e1C/R05jER5tyLcyoZOaUbBDreoes3Ev+hCWf7c5tpmzg9md1me
efvzM8JjzAbU5tFEir2tVCJoA2NrCUpzCqjkuVtXlcSkFa5tD++G0eAKuJRiPbQ+
bDPQ21NWmvRu5V0La30eawZqnPHQfrSKK0bOn8h/OeEuH9HF7umf4/Kb5Mg3pLwW
M9i0CEo/7Y/QhtJ2mRk7tt5EBNo2sYCgZ9dwtcE1alL9XGsMtn1zjRS1ktSsuach
+BWh+2D4OJJFJbEjwqIAe3vokHlmuTkgt7wtqqaiFunnC1e5OmwQgYZYho6yDJyj
99JLlYsSeH4AK1EkS70foY//o791wi1EuJLjXRIY6Rj8psB05Ih4VDF5pvOAl/S1
I7FQP/fNKaIQa5yoVPVYwPoxskg+c9M9ZqaxhGyWlMiIvk1TDuLpuMCyOQbwGAve
9erwRLjuqgr5t4hTOh2day7tqkRDfa7J9CpkQ8DICdL0bmniuQRyEdwhwfphS2qU
OLaHXMtN2+5EaIYdBA0PLxn6DebsRIgfFQLA9WFkmZuE6Jb+xK4Irfys+SsU5KOO
yBb6fiTxcjIAl9VY9+3P0jQwiebGQjt+/pcUFX6AU+7eRzyYxqNL8tcYyV20hvCu
qmMVg2cRtUI4KQNkLBMQVVDVFgSqvGe8BeSTZKPw0TJnY/see8TskV9+Jsju1Xc5
pgf4hwPLLSohSC0WrAOCWEEx4NkWCbxFw8Mdh90RTf6dbJv20WlqOOo8U6YnmQ1G
4R1UR+PXbz2uq8pfRywzoHXzLHceecfO/MaKx3KS0mMattTC2n3xOqvOuLFzhwoS
SixviF/WRXHIN5/2bwYsXnSGabNXUoNtQzr+QPpYMJ42N5DpEcL8Dv8jVE9/vH/u
CXmFc2+bvpspJZXSUuGeyoDxjXELULn3/+29bjL8xnuK4cPQ6vY8lsBo+T2OhA4d
csFYcr4lzwxewX0ZnRJe0MVuwJRtzwVCexdCScVbk9cAWoQzsqtLGBro0CZ0/+5e
Lbs7mGt0UdTvCOjBWZkko4pe+b4N73S4OfDt4i4YQectEpG501aGgCDPX5+myad9
Q0oApQcieVFHjx9yqd1d/s3ot7VGud9erMxbT9kXpy4mC5Vif4oehDMZgWx/qZGP
HCGKxnAQZg3DmHn5wJ+rPEsemCuMjtrVXJp/fYqumEAEaDR+FGiHxsEhRXXL/ZEz
H6xOfekelNBRZW7sGui0+viM9fH01M5dO+F3Hcz2bhNjseaZrpY+7vyU41Ow6jNI
cvsH8OB1wZrC4KpSrb676uBs9bq6CD/yV9cy3DpIMpJfVtEq2wQ6jpSO1FXI1Tv0
Yp6igMZ/a2m5/94fjHW59iaO/kV8NAgBzI6/s5F3WXX3kuIcI3zE3urQT+c7gt9g
es/AUfdKeNXfMqJz84S7vO6GThOPO/XyaHm3s/3dhqJOd2QQQ+++jgo7aSAM2Qac
w2ndLMrcDUDIL1vG0GRx/D4O7ErLp5z4H4xFCIyQ96+pXj5OeXO2HQyI+ay79tdI
iroLk55iK1UtyDoFSQQA+Nb+5z9bMvUJSnTHiWkJV63XqqhoZLCYGX/ii9uIq3lY
ByF7MjIyHP9Nze8i6TBLYABn8hrDhXNLmyiuiuYaUCGE7b7Vi/mQlPrivesl91v6
TwHy4PLJqnI/dTmiQ/uVmaDnozgkDozzMsUF9Hl/xotbwjG/rPkFIN9LxFlYnCpz
4BIr1m1HWzWxrj9WwO7oexaUWgqEtjtGW9b58b+KuK9FmqTCfeYtalVJrrrXIqGQ
Kl0KWoS3+MQycUBoORf99yBViP4Nv18xvl0VkCbNr7aO7UVZkDyobJ0TbFN28NzK
G4G6F+E/AGhXEv1pdOqzlNiBDj1Q6z3PCQIk6uObDVlTQPfwzPeyUGC3yAJYJpYD
GtqvktktMs+w1ux3/K6SRDOqc5htZT2m4cyYdBsjvYoPRRW5GoiZI+wt9MIyy+q0
dis7K+QNDRR9mRTtaM2c/vQ6RNTmK7lJYFbOOKGR0pVvs2P9HkOrpu9aekCGQK61
vcH1ceMGGjwEi/5hUhl34yGNbUizNw8lE1Lw6iiFSy9YugwvadsPZOoGbCOAxOsL
Rgb7OHRMq9uG6PHwdOkvDEjHEPi/2rWmkPXvT+cxeX9emr1qrT6gcCuxqC49OP4F
l4XvIAA6KshfuiTIaCHGNGRmpWVwpJEKOu1CEQlVZej7oNn1fON1nAM9YHJN+s4r
XOmMF3QFOoaw0A3Rc89X4fWXaOA9JHP8BDnmaTd5hjVD6Bm0SFYm6V+a5PefwEIp
eiS0kNvdKK9VRyCfYfV+e0f7io652hC7AuY+dru7N3g6ve41bVwkvuW5/SmGPMOa
RMrGhzVIPP5YWUtptQhDrqWmxCQXHW8PQgbWhIs+S+fP2tFIkhbwZeTGaKXXNQwr
PLo1l/jBq6FHY/M2rxmfhfCbhgPOtPr5G3/XAfyztmAIeyynjE5UIN2DJo6D7F0X
MdFYDP2Kvp7/KljviF/vArFZ7CLHH3GBAoBJKwR5vlqGRXeEfKM5LVxMHEev6V6M
9V3N+ujtPtX0FiVMxDST9ZF6jPNI4HBKc83b30ywRl/AYdPVQ0wqJHnkL6i0Z5N4
Tp6YgmIgs/AjIxYZPgoiP7tDoRXlzdJqbh9KrUb+nX66ALYLsuND4qoxwbkBCx+4
s8jwcTcSn5hxI5kJPunFDIH3zSRaWa3hdz3D7r/jFhvJwzhOurJ6S0qddO5Kg+1B
ZcLU4qSZhdEj4bJxJHc3BmZ+fOAYo5zPuE400w4TgctaRVIxDmP3MNheSZud/Iav
smxoOYlpq6u0cabLtrw0/b9SujDcVa2erTln34i5Q01oc7QrH+6A5fndjE94eGFH
iIlDsUwn0aZWS6rLx/O6cJA+206tDCN5diQ6Mjz1c+N8M2MXSLewoteKShAUEIiQ
52j/N5UezJ0ahttZOLTYhvZNsv5ZJaI8hXG8LtsLvPUDYo1kUTVdpwlpSZXhCjm9
ANGkpDafAImkLLLUbtONz6yCWPKXHV8Lo5OFFWQnBY8jW6B5DPEpZ3Ot5iTYxdYg
NR+9JdZbFf8S2y2N3+guN0sIm/wjy9RZL/n7jsW9PUWzWJShoDo4F+Qguc+ipPFq
u8nXpOpNlFqylIV6CvIhf0mUo+qE5H8EhAlnDi4iCYtsIiHkddp57PrnE7P2UoaJ
s8fZfnKA6PSr6ouLqt9VQYQ60WG45rYzv3TjQ0iTMi+1Tc605TLewCOb3RjCw9f6
gDFhXJd/q267KqreMX94JeJj2kK6gUiuKeaKu73jiqfp7qbuD+ypNtdVkW3bce8X
x9+sI0lDIxgrxbQcawrYQmw76uCNtg/3Ki6QGSoIe4v6ehILlVfl9okXAUqBzlSL
ntC6vqY+Sky6FlHjCQ/9N1c/jrquALAMEtk0timJ1SAj3ii8PUKHye3lxsdHVDky
3K2qpKHomrnG7lRFz/+7iJ/2i8LZmHtDOWm34DyvIeJatgE+kdR7fNsoDgXT7CvD
cZJwI6vpEWx01Cs4/4Hua7KTwv8QXetQOlCwvVJjPWFHf4/YQCWgIQaydchKHqYO
79JzjL1KsfqhocVNTJAfLZATdw0VhOZiHYsOHPT6YTiXpLOaA+JJV9hzD6lC0Vzw
1fJONsGP5tm5ma9iZqUq42NdzgnnFvUZppANSlfSrdG0A0VqUpgPQTjVShdKxT63
/QSUHo+y0Ugl7w6Y2UfGN8fKqV8a0GCp+rXQOS6+l7opvWZskRlnaKC+uGHa0avF
BfY65P2dSlbrZzha6B0yfBuSTPivu7ei56MPhupz9VWtCY3ZjJe6F+Gj+dsxJyXm
tJIvMID+V2EzPX5khIaYt2Ax/n+CgWlwlW4vAM4R87j7C6+p6+Bm3Dp14PKHkKrL
hhBllNyAx0s9F6lBzd47txIGMzleBfEOBLDo4aPxNhkwRNE04/Q6xATm2sSeAoap
C5NiAzEWPoHW7n91q+LSle0KuLMrK1gcGBuognQYgjYD/7IJhqUpyCo8jwG+WmZu
8Dze7YpYxNhrrtc+CfDYTzcIc4TAwzinWK3RS0weX9QhbLB80ghHaMGCh4X9kHm0
uhqu3nd6yENUpDkmuAjGV4nFNUplvnKi0QLKeBjiuJJcugQucxGYiPoyXDQcXfy9
LfYGphRZHdHP5RqFHP1/2ROpNNZHW9vm0IoOJM9sFqT4BGEE+DNcqZudPoDVPe6y
7kX808ypzcquwE8gHSSgJeDR/21gfijOBomb8IkPfYGFUAWyuz2lqEdQs3BHMCEY
8ZpxJtO0QpiMXHTwgmXsTaLUONiCHAz/qD23YvJiwt/KxmaU7Qme3LHWJQFsHZ4l
7aAUMaQrHul4/ofkyfg01EAzCU33jiFjQ2Rz5Z+W9A5Ba5y2tFTI+19XZ92I6giB
D/HIKkBlTam2fMDlAfUkN9t5o6hAJMV/wARWSmyUrD0WErLE58Fng77KbB3X2Bfp
X7q7l85TCSxbmyeQ397U+DqjaIBcZI6Jee7I7iBAPa/4qWYEOZfCuzuErDDg0B9N
XY0QGS+Ate3qPOKN1O5kzhF897RqGC0L3SvAWyMM/uE7sCyAOWCJ3kOIfZ/LPHmr
uBoBC1HdFYe1ZpPNp7XOEoAOXOEO5269AgqwH7rtnpss2fose8t3YH/ICgDv54Uo
c20OFUtxcqu/Uy8NMSKluXnTMwD6M+5y2/Zp5E3qhOnS0sRAgO8NEfSWrZi8yYl4
zALEGnF+bOWKtH7++rZNcefhB8pxdJyWYnjwfqm0ZNUa9ezjB52wtdER5QMCFJXj
yoHfpSEOToHof9l/XGUdNCHa+zx0X4UUHJ2GkGRTKCIP44W6M/t2nWBrOifObs4f
FE4f1nFX90/ioRN6KVHyqo3c1VjJtl0gzGwlYrALMdX648nVVGG3jp+f7yBKfp0l
QfT5uh1L8oACawR5NlqStByfQLIRvq1Ancvf/NCNPm6fGS4kJllPsDWMyXyB8oGb
LbLyOxx/qcT7zBsODuMN7Be5mnMBM4jtkQgyb+XuGz7+3kFUWwnWc7ZIEJJ4tXVE
fau05ZC0bY52nBwN1N4SLu1I25hLrnGX1faYKDwai+eYWya1mHLRk7lJWc6iy3lY
lcHG1BTYydbD7WQh0R2o+dm9w+patGrrJZXGHOJlHMtiNIi4hwFfVpvuWRZiLbpl
PCniQMG8RhC+0r6ZbHMvzdvCp3FuSeKipaz3m/L4T1LdeRlsubuVwdYLWAultwab
GXCvYRb7+xzwbup0qzAg4Gm+2fWdZV8P17pLRgucrZWj9HjtwG3k/VNxcIlCic8U
fVygAuCi0wA4eFPBHETFLH4NdMR7UFGhCSdM+pBDK/vAcX+t9HlQ4OEEvgsUzTd5
FnEHdjHNi4wc+8DIrpUogZWVpaHoxDJOjLTqcZfcN89RN12JNjTb0CSe3TGUr9FE
0LYzhv2nLWYWD1x35AnPRKzhtBoeyzcFhU3sOiSa+s43IDLj2vpYWtzwuRST+NcI
VPuKPcnrUSmw+nAGmK3amuhD/BTVuEORc4Mv0KNmxKDUCAZbxetDFhBoDNy+sfC9
ScB7PWBpzPjdyzLTlzv1qmIjj4H/ri0niWHX24u11S6mKRQ7eTAOTLXHkldUVJrn
kOm4k7DC/FGK/e7L+u1UwagQYrU31nk8vwfkXsP0xGi3IIhdPkCd2aEX5ETGcrEf
okEXt4qhboxidQwUdyZ8MW5ja7zYypVLBvevqzuauMe7e3DLznFS8fTcSo7OjI3V
ZaWLWluzbsDccCZGqp1US87PDRRRefPbolYd4fGouhdXUJxZEJCg22FPpn/N4dP5
41JYDdrB8SCXCWuWWzNVNA0SeV64pm2wWPDjEY/aiRYIbTrb4JosV4Hk+pIrEskj
cGR8YoEDWY+JXIYuXViMhpmpIeoU/NAvL8xkvpj4moQ5rglohWwPWVjAsMBNWA+p
b7rgTQIlfOPpIt/+fN+lvMjDZP6cRFCG0Ujf9CRvJXk0qVM7IaDNmKaWBFuCCRLv
32w7XOOmnnM9VkRHFJHZ7aS6LuJrPetlplQN1megOLsEisOGJdO7iHbnbFZGGSD6
U5rN2xeQTZXMktZ1MTZYtEpuHwYRz/6cxERByxgHtzXZM6YN/EE0XnJ/z0w0tZ7+
tGcSnJ4JZXvDCf8ZlHI1g3EIjnk0fl6YgQMjI6JmmcwNOe25Oq7apclMdoejSho0
4uqAf5lAqW7rshmq5PpV78cLSeOAV0GDzIW31ZsY5ADc8vRGQbnWyYAxxVWdXQeI
P7N0GihC2ebpZ0zuvTNpHJ4hyefccaiQlKvnvLtyfgpTmnUCH2cIKlwciNzEpdgp
pYqB4wuKr0i1+RcSQ+w3At0M/a+Y1xba7IwXKYbKp1eg/pVIjLmhhARnfzngBNqv
wtyMY3TgiEgRXgdl0meFqQ/x9C1QUsayx/nMmZ/TOGaYXgTaq+om4N0eSRIte6YK
6FE8V2EQCXD2TY6mEjK/uf/zB6lkZoFEqYaxrdbpJM7kIoVRkbzGr6ePhETCqDSr
WDxsa8QnWQ4gpI1ikLag7V5yzswKgITeEdAcdryMe4G5p7/HKEuXP5FA/Xx2A6DQ
YT1zusbK7usbkjfSxWLguJpTvIE0ffQZeVtpbkmf/4nJBvlX9LrOXjU+edeLrOJR
jcjwehw1QALkQ5LGWkkWvDjCybGqnirEFXCqDd53K0kS+pRogWVMrsoo2iiwI+F5
2Ae3C8eL1zYubFGtXS5yBCtGMIZYkgXYfIKnHfGIJvAqmCpMXK7VB/+Qnv6aF86M
6M6t3tJvpVRxvDNaAzQ9rnWAuUigWPRFCASpRg8+R6qA7WKUnCZEVUlfG5JOkco0
kTu/FSSGfZKYQPFr+6Jpw6+5t72+09Ye7P7HY8i4pVu1xGGhzCVHY0QyCBC7UW+Y
7p/bMQ+FC7oQkIranUSQUDs1YGd0x9VtH0Jl39NJI+L0SQeSlEYQYwsyy5warAH2
BjVE5MNhvbK/sQVTtAiH1WWYpZugweF6ImlT4W6TvLZuoh2zAcgCF1HOTeBsYsAd
ZQaDK2FtAEVe/cSF5xMpVoaYyTT/wUv3b/yYKymxAWbAqXvGXDOCFw+Zihs986VO
e9vOOQxrsxbKJWSmL30fW+YgzwDShdoQzBlOHCioxegJqhx/4Viu+NnB249DFQ84
ZmhXrsPhVY+7rwiSqOS45iQiCEMdlCe3jNoMeGY3Ioltj2a04kBo6gT9NB9icSEU
OHL66wUtPyFu4qVrDTPv4UTQaBIbkkuXbOW0ZXDkPvOUKRIopT5mS2nyaXLUad2g
0qN93V4bekpvogxNT1DN1jQAmAlZ4gp90+IyieJVQ3dgCdSXiyqrnFwkx0/OaUQs
EDXXQOK1ChfiVtin4sJkW0qS6xGmTpzVTo6+8r6JXQpJPvaaDCCf4xxlHhwRRxQF
59qYmHRABRsI6+ujNRWrlXysbihquk/Qd+GebOvySpEUuVBPVXecIYIL6ROA5HB5
hsq9hDS4Dle8Lw+cJ5WMowrzXAZDKFDHTRwAkuQTABrnsBNE+Mi4+zKHEUGi8u9f
42/a1WmvuZH/UsswyUNHjuVykII3QioexecSWSAftQOTgq0hmDQrry37CpleWUAG
Ybx3O1jcP2X9vV4u8bkmbCJypSQxyMcSDb7h5wSPdpyJezLRv4pmcTPubWukf+pj
AzLs+ccxFmUlrZmGv84Y7Cbh580v2gO4Qh6I0YdYiduKerJPM7mqBeFctMFh0jQx
3ibT2do+hJTiO21/HKX2XDVN9d1EcIug0AjoRkiovojUwi+9/L20sjwLcg5xxG7I
63EGkr/JLiPMPtxw2E9v0tFheX/fLEfP7sx+FHO1wuZhyzMmLhWyjX0JB7qgZVvX
81Lei2TpW3G/3TxOtfH2njDP1eQ/uMUruSc2EwRD61JTh5tF31NDBspTcFkNRAhi
AZoILXc15vPgjxKXfUV5xh6gGmgoRN3nSghAzm0Xn2og/x82qW4zLI6OwU3UOS6v
7okwQng5vQ70Y4RPLGD95QxyNiD90vkiQ1qLW2lVu5FJtTcrTTxh1n3ehYvvTXY4
I4TRARNDgsHr2y9ikE293u54rdbi7vRf45S/lq0c74om0N2w9IpM955pHTNRR1VZ
MI8Ouoyyu2EC+QUKrEdi5C3F5yBhfaPW71c0OGlXsb5G0orMXcDZSJGx427S6oo3
QjBSPL//I+Gq7aOtj888OZxPO8XAkwEgS5CGbthQeKHpK2uOr9W4bkLx5zBMUJ5M
isrCFOOew62Q1aHwUDmSUeWeX2hROoxuzEG4tzKHDTBqp2ZxSHBEfTGAReX+EEgZ
N5yaRIbiU7SIjaGoZW7Fig==
`pragma protect end_protected
