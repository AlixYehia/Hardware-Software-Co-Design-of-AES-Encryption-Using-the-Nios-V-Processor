`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VXnutzaIfJDVqCWfAv/Pdgd+6l9G005VI3U5E+logJkWtFP/i1LVm/lO/Ysl976P
8b60+XwzVY6BWH2tit+M8/WRUa8Dfw3AwOyFhslkf+HrT8+JXJvH1A7nlTNUHE28
g149GVsrAkFu1hn77GoUxcoxFrGwiJAKNwB8gZNd3G0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12448)
BRDvL8g6LIfnDUqx2WL7GeaVDPexqEt+5Qdt61oylP8BTZzP+vQBiQjz+f0UqpdU
5gD7ar45VkTpxRc9LXpNPrgHXjXBomC4qH1clfc6rEbkphgcgG48tEwsKlB8PMOi
DC7fFrWl2qjeWVpVAD35aIpDUguEEKU7AggBS9kXlve26Y20aALhba7D5seZ7kgi
HnqDYQE55zakf9WBnlCqSHmM3KmM07l6CgNkBM5mLk0NSfOaNk/xZo2Cs0Fuy7jH
b1lLYSDxMXXahi5T4+HNwy61am03Sz+trZu6OzB3s+hSRiPyc9lgcbGy0gmr9dEP
ICy4tNFiMq5J83+nORi3tZXIziZrSpzD7CWRh7dTf0EBiXFQsykIKNzbSWRFglhC
aLOyaMQNxJ8C42629PWVO1dQmI8Wk0XoldU8/91+JW+g/vAftSunxIvvqLUvPN+m
0dVWdSmBt2KBbhnpuItJox2sydaRqghZxPhThY3Whug9G9I9bHfteoKMhfKCn+R6
NW9tDwHkQcsvcKhpyVv4ExPWbWj5RhmipW++DnEn1InfQHiJ70RCFDnrXLp6j9WN
+mV2XuU3IexeV9WUgQ+sr3QTGDqkd7CSlNT6yKK+E4KKw6o1TQqkt1TutVfltGnj
E4Wj1cYJf8gXet9R+AzRPLCl/iHq+8JIq/bKxyG5MrfMhn54VSv6UiFHYXwq6RrG
DQuxwXqO0t98rphVmQn3gjHgHectLYE4bfzucsG+4GLpxF9lqn38/jqtPVgOqXoH
EMe0lJBIDgE47VZ+NnaG7uJ9I8M+lFGIrkim48G7owpeL1y77T32nnOauTqt/mo4
qudKhBg/OEJmR0ctUX9M1gTou7aAEX3jmj/g4XgO48eNz4IFT9MYuOOGRfK/JPR3
5ok9mu6CreM4POZKiTGm2+KBl7b4jYdOZav9br40S9uYPLOgaCxizDVSg2zdAX8K
s0EayPqFKbKW+w4cPbVZBDuRzja8/KUxUhqmO9d63OGWreK1EXl0T9Fa6KSQTC+/
TxgykAM7BCqQlLsaT2Xo6Cxn8dNSlnVkrrOvFHCGoYi8u8cxsAkM9MWe0IlKUSvE
iAB2bFxy3P65QbGzrsk7G85dDeNTqZrj6gUild/48ur9AWo1VMqkC/Pb4aiocOjW
4xSfi5Kad7fdzYBm10F4q4W/IPDXLQW7qJ14v6e/NY7G2zgDUsMicQdY2+AGu1Ov
/z4/RSNAWdsYxuZuyRrZbn8uWqOUp/kXIL3exZ0ClrsDTeTG7nfTfo6cUslCHUqv
t5vZu0YrYe3DluiXa6at2au7JOmTHztpQimHNqc0i/xjDuyjKrkPtEtklVvTi2K8
7RD7NknsyFOxR8zLeBfvqgD5ypUOPH5u8YfxeavXc7OzXCCXPWxlT2SRO4B8b3Y7
HUYF2f2wV2dPc06EpYE93qO+/TDF/opJHfsm56roL4E2DGRoYlfduVhezYOw3QKY
/EL09sWMV4RzMpM6bmbTgGkVLm5f/eU9Pngf4gB/gCZ/7hhkCrPZf7bk2enz7ieS
eHW2bd6otwjK2XOyBQhLHR0yI+d7e5gQNiDKBUtyTFpz2ok8bsbvjQtC3jn+hE2g
yYacRieuwjjl96YyAyJNbSAgJnvOj+bNBnEtC9X0D1HGFsbEjomoThvVNCqa6WLm
D11GFnD20/f5IICQ9Z/PRlec4UGxisFvwwYJj9GKqL9KYdN5U2xE6IRBF5OSZ3cU
LAYfs53wRiCmIZz6XkfDZsbPzLnL1TP1Vuylr/sNPX0X7R+1/KRQfFI/sxAT58vL
P+qRb+f3vUFXIqeT9KKIKZnqmlkWlrsZR9qQBejlE3EkJNmSeanT9M3nrfzA/V+l
8LDLCeKBvgL+qHYdMvATB/momOJnWdSv5YWeWGLIbYBwzMwWWu6EwEOBFqNM1wKO
O8yETzKrZ+6SruQmcah3fNMgpbqJ/Q33CAU3LiDMdfjDZW3am6U3s1bs95XmI/RE
iPMtFtgsn4QuSkoS0S3bnyBv6G2lTJSXAikhL1+q/qvI1zTtewp6+4b4i/JXJkEg
mxbSQtkws2F5MhUVhmQ/Zq3BrVSckjMadilO7aCcPEL1zjzJVaOGaJpUOmGHezFR
JQlvX8+4yDxR1QNRHSASUldFmrn8lBSR2ePBXBvbutqHuAr4Zn/4XmZUOBB2L2sX
RoZdqaKNnia8GT3QjvO/cEmTg0aBFk9wUawjP5I4+Yl/APMOMSHzPzSzdCEq3R/Q
96xAPeHOEPppJyh8bcFSKsLirY0Qa8w/4WFM+3vZNFU7rard6HQFTIwhcjaxzgY/
IUtenLTWyT3yFTNX4Tau6XPly9T6QMMeMlifwTGqYjBdvzXC8V8gzcYngkYDmY+q
vaAG90nxmVocp5EcbY1S109VvB9C617HuP7H3vEenZGT8TZgZBT8RqpDaO/l1ZkM
dfcgeDMTiBSw9jj9rr1vF9DWI6M1NtQlqi1hJQEM3sEJuoCtQZCZc5vSX5sbNqVE
rNKnkRNi0uXcRe9atNQfdLcIsvlNcm/6v2yaEAOYeJ3EqqvXV9KqouN/qD9xBtXc
pCgBfMbBX+XSmKOBp5z3jGw+K2o2Xkzvx7J/OnI9qljjFB1Pw+O6PBLMoloo8mor
3/oqcm1J2LnQ4SDjVvsVmu5IL3PraEdSsqgzDMeHzZd6vhEZAylcSMkJcVXbK70y
27Tds2lBgMQABtYvG1zTkBh2nAJJnB6wHZuPqEDLpN6Qal3XyxSuD291bu30LCYC
NL8N5Z7cOb/+ZkO4NZUrEtHx/+EHBm0YBAfLectUWEofuKT4rjwGcP/4VlZRMtXh
l1xWAgA6FAKKCC/TXrWOyi9+ahj+/Kbd4yt+QqlchD3q/7OdYI5xAL5SyL/nvfn1
blXzD2cUHf639RlNzkcP8F94hKIQ8DUidq7QlOKJUF5Z5p7vFQIHZ2d29oHx+cL8
M9iQM4i5B7wQMvxUXbr4uzcrI5jK5YH3/A6mSjgeQVOS8ys08wMqHL63r9ya2LnL
Z/JcoltAqMkrN0TA0U9YQ3z1LXZHOXx8PA87m7QihZtQ5Hm1bnYGEDfFt8oK1eSu
0CgZlOoHaLLPEP9Xlh6SikkQW9VBMzI+GPKcjwwVUQyuJ/fU+gxu32U7Jqugtzd8
BS+a+sFgLAHVR8C6Xge/s3BdHzkFW30i9aqgMcOW7R8wZmDbnYz5o7/pDzpJ/h6r
Dyolh28DXGMqI3cbH7UNAQsBeaseIPOuLka8Y1C0vYeAIlytkIIcJioesGfd8cbv
b+vwkAu4+QrMFkysJ1kMrHBg2+8zyHWfiwXXqWjwJHogbDadBeUh5xdq4fhwQcsg
XNqSjnq8mnzgRCx2tnB8RPBBkfittSFwz4b73ScXmGz/eLdeqLGzBEoyDbKiMBv2
KIFz5rnhKh+c3+RzWAwm+VV/gkOR9Lb2PbIk17Sx7TUEcCU/+vD3a7i4DmPRrQyY
rorwKgBKRw2/s5s2Do8gxzR3jY3YIr1YxViyVsGyFKwdoib6Vc/a57MLqXBHG+Le
2deY+44nIExBCGuoM80VoCcd8BDxV3sbBG+/y5p+8hfxjaWIpP9LmEvoOG7vF1CU
4c8k+OcmoA4fzhKXmRLOiYm9iFK7SuqSMvEOnzGhxFV/L/TpnElOLszN/Ss6k1+L
9L8Z2MKA8fCl95SoXSxyLr8Xc+7Hcr2pLC4XAOt+GdQsm6ZGsinyeU78MOzHHEhb
BeFyUfrwbDtGGJnBVeWfeURTE1FpIMPpHG2TdCIh4rT00XSdwmnPREW3VZwMLYL6
VjnXAJCy17QhO/3h+E8oTPlJxLqYySUKMcX9MKJvFNAf7kQ4lJIzq2Y+DgEZg6OF
cifMuo1Kmhy8f9Ufr+PtFJn1kn62ny7EFujyfT1md7MtxBTdKohDVXWvutms2z07
UmhUx4QsyWdnx2n7iXVAQn3k15O2BXly7aE0bRAszIMP5BJzdMJ1WAS80LweiizL
nqcGK6q1jtscPgf5N1bsdA++NDqhgXgUNkQJNDyaS6xDq4FyintFGKJC9CKQcxau
miuEZh9pxt0z3GnA6qnILqEAXB678gf+ER+BD1ObJ0W9cxGWpbx5MLCKoQ49szh1
gkcvwvzvNTe69+dZN+oC1AlS/JHB/xLJOvsR7w5H8eMF+BRcTFKwUl8vJbnZriB3
RJKoZDvk4hlUZtC5arGns7VqMgx2+GpiuG/OrZMn2Xbo4FLFRPa8fCqyabV0w9xB
MSeBcZCHR4F1D8Ug6dYDc4RwdRepBsWJVgND1C0jnJwlGEh7BQ3ou54b2nAWAf6C
EpEABX7x7afiy9vXD4LyWyp+H8t4FrlbtFAukPMCBMLPfSp3ig6PCI8ptQT8qNCn
Ber2QVd7ViIuVNA8F7m9DitjLDmjtodJztvlAQ/zqwlUqRvMd6OsAdDwQ+11ZNOf
4+okGJnf31kkseSRD+vOHs2mg7eg2B0eJy6eWgJ8189xtZY0nBkmksk0fek3yfUw
IBPq08wh+lBgTHPMCsmclPJuxCNCmq7UiqJFjxK5DlM0Rqsr9HGRIYZKD3EIoHkD
fwV0+DA5Q5yRCbGK2LzBmNIpQ8bhS8b+cJDUsJgGTI+s+i5N0qT/e/ARn6QHEFX5
zWkqocSqwRCa9CTggDyCcydbZMddpfF+pTPTuS48LA9ahfSkdZjUvfXbUEDhyBET
b8dftCnPWm/eAByTZYkEFv97dSZ4hUfEsecE5qFcg+nFyjjtrctlgFWKl7j4vjMy
SmdNEszkGH+srhWy/GTjZ8a/P5fttb1lRmpPmpgg3d1r+5s/0Ptsfg92emlslLAD
CAAHdQNMqlbc/nqSsc0adKwzj16bC4gXwQwRMeAAzTGhZWhUHaY7MtSKbhWk8Bn/
JYw4jPO72j8czDgOUZJlrsLHLmx30dL549YlDpuKaV8ojoSWo8BawwyIIfyQvyf1
sWdyRe5BNpdGKoya37uFYPeoQ7y0PXcUsWeeGHV5+QUVXhMx727wzUP73fxUHXVY
Q32Sy+iBjh29UzzLQQBRiukFrqOsA4UHXaMMryBijAcIpnU+jeiFjXmbMPgo83Z5
tManmrkzS4wPDKQDSxWBgAacJOmtcyWeS/rmm30973ERF48yLZtRU9tR4ALNEdw7
Q+VQ5VSo/PsgJGEe8O+Sa3gbl8bjdWhCVJVqSHkqV3sbt1B1/WyAl5EZIB+vf4Rc
m9jmOdfRHWUCSxhhzv5uHvT/xnBpZxTw3bbYDHyQGkwYAEyM8ngzbrf/IWipRcW4
eVn1/MG2inVbYNyUOKkIMp+hYKO/0eQDFQ1QFpn1xCsQbRSiCcOvX4MPre0XkGj+
h7Xm6j3OHg8goe+brezbSbNZUUDboryDTPysbmQVOsYsZdCH7j+OQ/zNMP8oWbeP
IbnX2xfzm9ooc8wVrtu+dMDUhTt63nTOjviEDqnyb9GjzNv+C1xNypYqb7mEuA+W
XlgPqlrcXwsvAOIATq7u1CqmQfcDbPTdyrjk54ZaD2dyAfJXJNNvYvrpQIisXj0/
u0D20/WGe/1/qDb1WpDsDtxmBSMrHuB2Tt5wHrdj+nYuGQitoylFYrPb3d+3zWz/
xZb5+O5dRZxAvSluMG8dg46myJLLrOIv9HodFGRA3aPywpFuwPrw2fV/yzJ2T/Oe
ZDfOkXgEDylQg95GNwzpuj1QX48GitNy5bhwNVa8QEoFw6OnRgLDGDaAnft0ojps
I5++Tav5jdwsbpoG+YB2KJZB3UTgQYjvd2AoJlVwQWw/4oHCvkDuaHHSXZjpDkK7
NmGsCjZUvufpwVt3i5Vb39LxRlzFWYanspFc6lz7JniuF4VFV+aie9aQkmZc9ID6
pQpLH1SYfljk3C5JOwPoWr8f7U5iOPjzIoMxc0DGBD2h5mUUbxiQYZOw4aBEy06c
+cK5I1RD7p8AuRp9XxorI3Z/oPtBQ/XxbE3ETg6jNQrNo8+5twteaXLoRl2lao9Q
ROa4qJAy07zUASGzu2hKnYlyDNuQ4NhRsMcLeyNwVNPszKjEiNZLyyBfdF5/k+jH
l9OHR5QQqfrJ6GzOm5y/nQesJ6IwJpmFLkjPAexccLLLL9aqu0usULCXMa/Z1dks
U5VDcFg5qhvFAbCDD0VYFSJPaN9DjMRAUBvC/YzJ+Qqtj81S0Q4ngmFp4uhqY4uS
xXw5XqSSLhYCrWk116r2KoSn5+ztPzBp+w220m1sA4XNL3bVniI5SyRRmZM4anzH
y80um31UtrrU9odORX6ac0unnCt185tebp7lTvtuHICe+uynY5Ha+YuGK6wzq2gW
gvNBYzybp3N8/6bkSJpCZH3kZLOpmbDfap/qO3xuY2bkZL7fdqxzfxBsbXu4VGTk
oEODequVE/5tPFLFPDpMXO0Sa0eUqOgyT10CeDKUZE/fCWOuYE3FQTQdUgcI1kCV
Tm3WAY7VPoOA9Qx+McPXB+uokjG/xyGHzZXMriSkhctNlqlmUVjH09yCnPjDoyMQ
28FTkjXbx1DC4Go6ic0fTVNY/h282ZWELDM0TWQxGCWtMkYX25EVaxPWAa10OuYd
fERh2wGGkupSbAfw5tiONGRA5qm5u5Hnq2MViSVUmJjWYWLRHuTmZy5BOB7xogdO
Yikrw04HeXpNA//5BSNeDn5+stP9eQhNfB6H4wvTUWEjr9vvviS/Kh6JaorjPuCT
d4sDwrSG1fjSfaPrlI/QfJdXIdQqC2Fi6jeTG8vXr/9D0/xg6C/jfV/05FrzgAWI
N1F1hX2OQOf2LzCO2PTcCgx3y7Mu4f3yj59tVOpgAa5yOAd8CTmXp70+6ma1FqAz
SoncFyhpj66tz54dbIF5lwzZHWa1JE27VAYMci2KTkJmS3Y9u4k6RrF+Rxkls2/K
yQTpP5m/JkV1UTAtHHGpf6cdKKJkNNyacoZkA/OOaREXSyIAeD7iuXyT3Rzf2S8a
fbjmEqcWYL0lwsiPAA67m5WsSCmT3IZjwQivckt0Dy5midGmPY+j/KPFD/gYTduB
8N3HjQHAAhtu/CdWrw6ne3Sp8rDK4TzsUqXUsvzUvRjYJ2dLF1bz8s+H3gdA7+Qe
d2inRDzhzebXYO4XE1PSBog00B/moM2E9dBxiyrrYPyBe06wRzBcCBDMUmx3GDLh
R8r8cgfVt2yC0vr2S3eNYqDiBOMNn66Wc+h3iMt19Sha6C7+HtUgltMyeJiHLbR2
GYRMZHi2mXb3Kfq/PVjtqFvjO/5wmE6jg82heSaMsWMPzZENadMalatbFFfVlwD1
0snNmr2hY5791hgJsDuEKVgWzXt8cN3z8FyzzwEAt5IYF/I45ffrEwP/7dEvaNHb
FBOdSyfxA5c9dbgcfbzpQsH3vR3olpFc5I7lUFI4ydQw+mP88RAOPUeU1NbrJxU/
9llG/dmVWOsw6MZKwh0fHGRwCVMAAI0i+JQnUNyBwtsLFVdf4jBhlNTtBpQ0uDBY
3rE5XpeSTXwl3cuWAjGg7ud1xGjdET11EhE6yu4sMFjw/3Tqru7kHMSd4gpNM7Pw
lMeWCvMMJLQJfOiyvQSH10gQV7v5PBS8Og5J4H6l+Lqx25ZOZ+P70yGCqp2LV2fE
FnYOLWVSEgeUWfqpDmrfvgQtZWjxTUsDikkrMsWy4RPjIusve/t7p78uaIVIRG7K
LyTlXCIRR/LENm4m7LNg0eG/jDQcumetuEazJDV0v/z2MO2WknqzJMT1qYuuwefI
H/su7lALUDyFgumdJIS61klf+Ek1ShChhp7UGF8HWiIZ16Bdaqm3Az/pgWdYVzJv
Uad5qyqH6f+ZVyMaXuHfE4onu9y+I3f+4aG5EYvNX+hSQSJFR8yvAZ07JojnVk+T
DlOl0NcuUKpPrdvuRGezcqT/01U01ySiAffAtzYWYJQBPLaVRVy1f7vVdlJtn2eK
Wwfw5AZr1WH3NK4nenRkWVFEcIZlhliKFccj2wBePzgG6kEP96CY8M6QmaZ5nc/3
fBhFYYNKwIvbKs150xaHkTPL1T9BNoYSgm3SZ5EGREfAs/EdkhFqQiixzbHZ8fDf
CNbo7dnl4JgtxW4nOQ2Zb+0U0OBS7W+MsAN6PmhgBk5sgf00WxjXizdOdkU9YmfF
Z/aP5722+yf9jMoNVVLAaTM4e+YrGiHFD3O42j0gofuh85Ugt2lhae4WEbiMbCYG
NSad4aC1N3YhXByTmoqT+RmQcN26EGyeCQeP4OlA2zX1XWyvvPI0MU5bylIQxs1n
GzoXRq8Ydc/nWtm2Wz9gzpMJvgBrvKBNNUoA3x/WqPtNG/5LHhg+LTSFKe44GpnJ
EOZZR9Z7mKtTK5vh4ONLMAN9TZ2wimivKS94CEnjKjuMFK8qSe91g9/wpSoLaecT
tjq349JBPkAx6y0TDubFHIepcMnr2vCF1wIhaXw9Qq2Udj36eeHX5XrQH/B+D9DN
jwWcFGrPi46Pfxqsi/GobM1Z3eYxwVDhLRtTtNJ0TvGa2z59WnsWy7EZbXpA2M+J
4RrwSSTl45y3eOYVGwlCTR1X3JoVIlbBbQPIrnBTOeqq5o38X6cEZ68gQOidRn3T
oXIKZ/okgR8ZmR7KyaN9EGi/CGqeAt2Avx6RvSR7YnEZZ0WyUairpA8FkavEDPRO
gxbzZseVap9dzJBmBSZVbmjvbe1H7OU9MxtcUh8xnwYNeQRW9im6+U8SUhNmvwJs
ax9ZdDdkeYox42GHjeUM4w1Jpy5KcUifjSgmih9Ew81JjOQ3eEq7B4iY6Nx0Cn7b
87GUisNIhdIOZm+z2EWmhRmWYD2GxpesxnZXXNMFkbul6g9ImRovzw78k8MdM/zO
Snj9FJbFqUKlzY0EDOmGuSs74um+AYC1Ejsue+6iEKhQw8AW9x58yFb2d0hQjN3T
D5TBcaXkiZRN13o3AuskBr6RKfq6j2ni3vmUORN/njCfHBgNK8Uw5L65FYx1ibUz
XZPNdjGPIVKJIWo0BI/dKTwf0SwDYqcAm5Bt0TpWechFqIbNJABqJbm/ewLF6MTL
QaFg+fwSZpnPRlfTcu0CEJSdnrf5CVftFhkH32I43kpgkH8x6787oAtsWtLbAM9G
8UzBzb16+3jLqsLo94b1h2xC3iYw0p7h3EbGdprr57cQZ6TCBmnLB4+ZzlPJDpwU
DfS8oTpL8t1sju7NOSGAZqdieu3wjrsN4rDdG9DsdWUvASXMsOMRjYX9HjdaD1Zz
gEhS+HO1zx+ispaGluczYJp5fupnGKNhp/4Np/XbrsV+pu02kXaeDv2kP8GpmfOP
RoA63rjydilucYJsCkwGIsQE1B+N/xnQk25w+WyNLEacug1gW4TWbYC+aTSlmZtm
igBpukaTOG1xAsmj4rGMqXzsAGV/wYVu5VQ3MWqlRMq8WFFezXeqJsF9l1TSgBKU
QHipCUDoWP/5F10To1Xb6mchU57Tms+gDo/ryzcFpEi5yTmavsdyq+NUp43YWLsE
3hApZatHv85sYBR0tDwYW67AQhCsEsU3e+A5tWKGLjYVhR/IB7KE11Z6wgzrDkkY
+Lcknidr2Te6hQHBxGZSsFUOTW3OoRXqS8FhCMG3kb7S2P1Kk59AJgcBT4MWjNtY
p1suSSTcH5NRE5WJvryHqtDCXB4i0sRG6+orsDZqWL64xd81E9m+TaTjM7vq1kS2
CgjOWvlXLo6sPvq3npnsA2NlxvZnOkAMjPBqQXepWD6ypZG1I9QKi/y1xq/lFxxQ
w3gvSL4PK7oweE9NchyC4gZkksQ85m3DSNb5xzgRhaEVtebSTuEeGFDqIHuLuOye
tH4xf85fuEiz150UggrhRNsZC6bSB+ClSR8BcgpMvgptUOefL1lNGVUd9jceWo0L
Da+e6plesEaJC/6RogNHAh7qWMjYUB0qpfIEMAb4oZBjcgik7gy2m2k0NLmL0nMT
KZXj+P6fND2AkbZdnWqYaRaNddgBImEVEHJGGVp1A3Ws088l8gJVHISc63+R1HCB
wuTtOk6Y0ARdda985TVheKg30R9bJnttepNlWvFJDk2H+ZDMSyNTdV2tr0bconfl
ICKJJbZ4HyniqKle1/Ga5sQLw64PWRKmftq3aD6KVrwU+D76BPNzmfoQ9xxkGCa2
4paxY+3fUososqx1PxV6tkAImovu8PIfwD60WalGr99n6ywIrrknwfnTX4RIy5nL
c0d4wU6DaJft8cngRPBtwGAVP5pGWpnIfWAeEI0rSADxYGt/JmJkqgOuVVwoUJ/c
tIIsV8OJPYywo5BZOO8mpQDUgsM89Q1oEK6X9yHBhASJ3V/fdmF7O/Prxx9aHF52
fQLZNrm4rqNciragFo5TY1RLPvuN2uwAdh9BtNqa7LbWK6C0iX/PyM5eCohCr9xU
ITlK4bILQ1n03NSIQqLqkyDRFkvZhsSndAefVetu19EmWXiVP5FX6AoNjaM56wxb
TXFoX02ZBylbZGNCT+JslcfJASwUkn/D0HAxaUN5xhKW9qihXVzemRcxdA41bf8P
I0k6jigV900dzmYLLPbRAVLQcDELUHSGgR6v1q2owu+GG8RDzZBA813hLXDxGcVy
D1Gntmd58PecOCI09YN6luTCxWnmVe/otxQoK6AQRy9RvkFEbVhK6BgkE6atv3Xm
IEUdU0EG7O7zCWWiTnv/u5RbizaaOzTTM64xk/9VUo+BEthtvL4EfC5KoPqZyaT8
wu16pr/NqgzqAl7PFmSuubkaja+dgC3Upe7ouveBGOkX6wFZ9Yi+QhWoPhnZqu/r
n/BmjgNl8p77nOUf7Qzij6Q/lGRRlDckZs4sLkloC1i1uSXNXd8ov6HuUuzFp5P0
DkkC/7htPLJVZGizNKd0uiNK9YimygnF8k0jX2hc2/LHn/LTZ+ClgLC8rlRH0JVw
ry9Bg+wSi/ryTk2TyDodeta7I/OESJ3g30xOFbBKkL9kJIlik0inFsfYm0F0h1T7
3hpB+jjZEmzSx9e/OJ5BQ9SBMbgfPvWflmPomUPpsYnIeJETZfXKAtrYpkDSBzjK
BZmuZ4mms9rQS9ncS+9qN9HKuBicfEE80tVX7ObTdRrwa6ymeYahTsk1OoAAZkeR
GY8WKSQvd9/2qBSqHOh2lCJr6HMdp9Oupc+9PPybE4G1BQK+phetPQLh1itfD7Mx
/EbazuPAmP7EKTxTUPSvoiJXucP8XUIUxz+DW3KccpWIPlziSkWOZdM/fTSY26tf
PiQnwdP6vz2wQi7Jd4WoEHyQ0PcG1Ijv9TgKXRkmupS1J+S1F5tel36gmA+7fcmx
HXxooG3F8org0om3WoQ5tdZC/aEiLuw7eMLR0DXgyD3gKy2UCKKwKjZADgMUQKJ1
IbrMlpTtLPPAjLLqcyxTykozHsAomOD1kAAS5rzOYublT+RL8iuYYuwFiV9BhFN/
9SDp/9WCXpa85JMg7QNxYqC79sY/u9/qxFLLj+Qul4sGmVLr9WVGsyK8oysfmXbP
VdxqqGs8BjI2X3H0HYmYTdMWQsINfDzOOaMfgKO7MuS975KonECMROCFZxC2R0U3
y7+YhcKptADMFpYEQJvtJFhfnILnfxSsLokoqQ0Lp7KlMZQ0dDRZw5EUlwpATzlT
GqfRexJ/TFQ99rOOh5RW3d+fwxt3Vw3B9Xit/lJuvjnhfx2BlZ5p5DcYcGUK3fT+
YlluHUzwcS+hCdfIrmcYcTdwh11KGPun/9dTKZW9FR0yhEUbWuwLlui95U0p/bu0
RDXqd4RK0TCbyYanbLItggHYNaiygA08X+Lg9wdXsKL/wRGyn8OrIvLQM2MWKJW5
PI6pyAxSmcA9j3BZoMDGPLn5U6smHTdjO9vutcP5Z75j7iSnZho9YFLkw8FKfFyE
XIWfi6vwMpoizDG5Nf8OBWhecTnZxYqWJ3DNQG3ne2OAraTjnppok20xPP1F8Zdw
Hw4YqbK4/JHWxUR8xYHq39ZoDe4mGhe6iKjr0fjMYe5KrVN60h033L1UdPrY6/7C
weFcTPeWt7shsmCjmQ4AhJKN5L5ZDm7HRB7oBDDR9RlaPZshrAU4WRx8XZdwp/x/
kCr8lfpWAwfoo3JWFIz1bFgTyv2DoSkPKX/PLRRm4u1Rw30u/EQ20zLuzl8cX3Xi
qfA4lOlW0DbHpbFAPyblgOHabX/yLaM3avKmrVYiqpr/jRRTEbnOG+DhzKAkqmBM
7JZYuYQ0XBL8QzE1o8f22xb7sbw8QrT4lYWeql2Gqmj7hddsLJ3lMrjBP77xqDV9
Cw8jxbL/68LDAgPbugCTgY+Xn3csyHLPWcjYt01WVSBQDONNDsuhk8qOgvzOoNGX
ZO0vHy83hGX4ECQeZQzKnXDV4iakgGgcmjZ7KXWMT/TSeAJnLxxdiUsZs3JqhSg7
hd8xgF28d2aQlPgh2560tLijUXgy6af2u4sgbDsJq/cp76iyAa8PZvYfqukvc2Qz
wf1l+LylEx2XFiUFQkI4p1J4mSWIUKeDN28HMiUzZbN+fW2IPFG/9Abh5WWk4kjg
B2OXU20hEGGAUeK2xXf2XZ+SUg9MKTd7TkeOS8ctbAgmLOAPJTCFIaV9xXdp4VJt
RdU7Qj6Jxo7VjMusNkuPHN60CfD8C08+cgCMQrFQxjRoivZs4oMwIlYs6AtX0/nJ
og3P9Bvi7G7JgBqUaCUn5gxU9SG+YqKi2iNewPv5LySrU5Lx+eHKGX6EOVNXNUlC
u7hyWcuRUJxHN2YwtUnq4IugNRI5ny8xUzD8iO4wCcH2Q9z4cRklN/qb8pi+Pmvd
GtHF8AovcgqBO4DZsmtUj+YbhzEH8ODTwF6gFnAm84MBz3fmaBhnuGr1pidl1lhR
crC87mTuDQN9y2KvMWiUNgAhfBBN5FPlncbwCnAjMsUOQkrx5TNUbEhVTjLGimwg
AuMYp4wEP3W15bhUbW7GnH0w+1SNdiYqizPUWQ+eZPCG9jPsckhhBfXpsaSJ0dMo
JS/E7T5Rzq2+nlcCBt0lpOmV4BfGuH+xeBf6VBM0AU18xgtQdGqKqR54zYLCC2Co
pB/2j96HreNnebAA/l8Majs8AYli72AowmugXH05LGFVMslWCF7JwOJrTpLf3zDR
bGyzYrCO3uRJ5vTVQQEyzIqKOtpQqq+wSSBR8tYF7vjze9tPtQhp1WHCHDN/Q5Nt
BZsAwe6jx9YYhxelCMr9zRQPtoUAm24bBnOaPPRxSP5ROQUkZJmt8PffWU5hwoAg
7H0C/zqAUjwV75wnFFMiOiggABgSqqQqTgRBmdXbssGo7SjZ+w01+dYXBRpHMRHi
4zq7lZM0GV5MrOtvfSqykkyOcpjBhXa8BPzSmmHUTCGJU+FoAcznfUzEFRA9Z3nS
eoyI0xC+8Y1ZB6zu1yeJtTSdGsGFtRHAg1K9hauY5E0t8Vm0bjJG16QeQSBQ6qvv
LPTuR3tWf0cBoyGLFpSbZrOsTPMOpZR3fRayv7fPkPw+T3QXAaUGV1PA8LIA/UXr
9JXANiqzVg3ALIsVGdohx3Z/TnLy58l+UyETBseqCx3nMN9MJEA5A6WMsAW9H2Wx
S+wiJT/Vz/TawUIiLyKiM62SYdqudBe8Ie94i2Rt8zyj2nU8ODsdxGaraEF0d9FC
XjYMmo0WkwTKxjWBYxq3Y4glZ4RpnwsK07StN+FVZyvLR8GZ0HkMZZH7Jwtr3OXq
5aLDiJUnCxv3wdLNKk8Ctg0a588QyBgsA2x6b6qJo+1xUq6SB1O7H81JzD3jwuFC
LcDCh3A5jwaX6cTiXv4pztAZnHdET8eZFCnwKRV/JdNiEJJcPB0GZlMqgTbX4PMk
c6pv1A6F6SCICeRBydegDj+o5AEOt3h6jOjFW0VerRSDclCnFTX73H29JAERQuFd
XZMchRMg+iL/BcoAXDlmoIoFRkmYuIc3UNNU80RK6Nb0nYwvzNQkH7MFbwBssZsT
rl0MXaMX1h+vox3L+1vp+PB3dwpQiWG8+9Kk9XhB+i22rhlVqpAWHQELFlTD+Qpq
qgoIO9wMg9pbXTD1jKWwFVycOmUuC1pYNrMp4eWLzYPo/1KSkoUc9Y0BhGXrhQFl
DwmckL3DpHdVuB3bpFX5sNyt2NyVwXpja9yAtPgG3X6YiJ5qwFulMjCES3qyzN8y
RysKo9uqK1DTG6XQjHVI3hMWjauhWhjs/higG87Y/p5Hoo9O0hi4lOKDX4sWHuxg
SL5XFpyJneUz/o6Kl71cRcawb7KDBF9vHxuyhliYdZqO5KzfLCD4DN3lodzyiWIF
M+MuoNhS4PiSD3OrNXm88+wKMm1t4E9kKrVKIz4TeSqU8z8VYZoV0UwtGem0RoyK
59AOFdMEYViWsbAx+wuV11tBc0vFRfK+SWKHJ4LW9BshglSgZsNRjC5nV0zeO3O9
FzXYh0U6bsifVTfQHxMQO5k7Ec/Wpn4fXhnmGqituoU850KBp9F1X3qme2184Xff
D2WV5RrtkusJyNK6X+YUe8giDBm8jLfe/ysDEQDnHQzh3DVPDOjtDOdiFxevaEy8
SUmW34b1pBg8MM4fEt/IqL8iFqgK5WYui3MS83HrvdMKImbsxvU2IStla5q6fxek
1czVKiwTS/G6aPJ0O19kOKOpvqX/b28IsSRvNWfoZTFZ/tl2f8xEIQxQcTzFEuaj
j6ShhJZQF4NWTS4dTPAiT7kryrBmN6ho9uD1zyreMglc8fjLdh1T5/K6PNhumSwg
mjyCkw6n5BzPlJqSDUby8Osm+VOCMTft+EXPnSVaFQx1SQkXATtlZ5r5KFsvUMgh
kyZbxlZBQ9DNdRYtDC6Z+XCgpUI6fzd5nyBCqKVhOtgQ2bGOuygZnq3UQ2kEjgJG
uIabQPwcfOXYw3vLQ9GsKmYkt/3EJ5i9GbzYm9PGv8FbNONda0Ad/9wtvs8Ag7Bz
O1CRdi+mk2LvSmHLbe1VshIjtM0fiOH0pCpYvP66V5IJ07uJIjniqn/cdieYAx1C
bejL4atnqbKKpJFuVco25u+4aIbUsmkllLd9eLP/nbhvLPC4HjE/q6Ea57B6Pc2/
3R0rJ1twGtmCQbQIvDtijtHikpCUjnfwbrhLGqLbiCwwmW3wjk/LJouhdZat5x0d
4m18S3vsdjNzMFl7M9XxAuxhWDSYVmUIlPUCenh+Hv807GzIy0aJz7G15XuvadtW
Dx+sxUwAh95CDhW6l2o6VBxotYFKJSCC5fjY97G+xOgHqsJsjy65PHa1fvLdfjOj
PkGxp1iyNUEVTNfNnQNo8lg3ubcYep5xkLLVT/EURZwbssfULJScF4Q2QyDNXlRg
ldqwHEAPaGYer68DbYOdSoGHwYlMmtC+eiH9Lmlw0oNCWnQnZz3a9Se8Sl3fiZ8g
vhJcFbIBEfUnf30yMRsjIVlvcXLyy/sDGIKpoJqFDpuQRlZ9kyXp+M5QT3+U92nE
1kNBBDPxjdQEqcn+TwYJJ1c0XNJ/rIpAsUpOmaqkekVPzu9U/Cs7qRrzfC4ZSnFp
qdoThEZj+g1gPeKeyPADLlpG+VIFSCXxPqpcPCivtehYMxa6Y8JSyhiuENcs/sRl
c/ByND2giudyyK3EYgfFi73vpYbLhX67Q7jPW8AHcsEHRrNiLQj3jp2yd2nlE9bu
2yFgQDJ9Oz9mnyDsoBCNbr3V0Qp5yqLxbTDrmvExZ3ubyN/huC/2DbmjWprBvxdA
NaFpiwh7X1I1DSTb2GKthEfj2mIcxaCqeR4oo47yHA6qmtnRkpapmZRiZe3VaHnK
I9IXl5NJBPCo/C/0xWC15RkJ8QxZ3JD1WPJskKRnqGL6DoboZrSk+T1KSXqAuIW3
8I4InG6xxzYdWuaze7dhuI6VriMRqhXukwVDodz83QUqoxBKnlL5u6G0rsZb0WFr
FUwDHT9V0ocFGyNvu0auOBAKpJ6ycJfn2Rl4xR6LHaV42D8d1GPxAELT0hCsGoQy
c1PW9RZuvKSokJyCJj2OuK/qq1lOrqmV6A2CdGKxEJHR3qmnsf5xGMMzKP7BKgcd
DKRCCSdAagEKnV8ShrV6X7/xTvG2iPeUPY1l30f9P4ZjOYGACvZUaOKbbqLrnICk
dRgEjt/uVIIQ1Z6S7ERbUMHDMNJbLy4w6SrDxUAtb3sq9tCjzAa/fofORtbHnZ+T
Qs9V/xtIS3ay5YSD6vRWUzpiapGlcYkAtBJ4ZVKdhTJVHIpkm+1qM8tkgyJWbBLf
Lg+IIhbmZjeSe35S/+0Txq3phIBydJ4oQbgsRYB+A8hOZHXmS+F6tFUIw1GmG55x
lQgeRjRsJYK+dsh0NX46kwffOzdD43dYaXVCMOer1FD+qdNz+QCVGj60e3jDVTIz
YEyRU2rVyP0C5BfZv6aZy0aZWOmOlD+RNt8bEEJOjoNMUROtYaSQtsBVvEilgq+s
IgM5dNiBH9c5MVQ4N2a10qNgTi71tAlMcUw+giRpjxa0K8iwRB0znwSKapGMIg8X
MWiVbArydel/jefGQbNm0CQaLIuqm3a8+xegZUaiJ3sEO8OfOPS/Jq5yUMD907yD
Uo5UEjjiW1HSdLYanDBHDlWyWzvmWppLzg21IDN2mPQzRb7byoobzv6Hqy5S6nk0
TutHDh7TXAYH7s1fFk9QqHudZNWPd6ilBiAY7bBvSA78XiBjrDq8MYV6LYkkaZvk
vs6pNw6cr6EG8ckvOgx+lqYd/CfeMBb162P7fzqw7K3LROU6QunAFJShnUFJncTh
OyXQ3X/6Wx4FBf2NQOVmoA==
`pragma protect end_protected
