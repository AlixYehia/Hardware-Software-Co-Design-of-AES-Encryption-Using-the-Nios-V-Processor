// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Rs7927gPBKDkJ3smLsMPioyEz9bLyxxLmoFMNxHg5HMbW5Zy2K4UnUZkgZCDZPfGGxQYv2p339Rh
QYKgA0q4F9Cbrz/Buc1d/SmHxiBZYlxc/ICz0ylBwuNztHdFOtpaMKG5azP1GZRE6cO6swQW4H0S
FKH7s/Mw5X7OQ6CKsCe4ImxeqwgEWRcZXLtBY57lsb2JBtyvRv3kZSt2JQNykAcDqqJrVwPtdtlW
mAb8xqdSjcnLVaQJkYjgxh+USEHBJFBVLGlmING9Apn4z5sitfO7O8AkjGo7NPkQej2+BPIz7PZY
9KmP06KtzXkh+yAzJ/lOzTS6iSzPAUc4yrj3/g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6896)
dj+/GtBuexv6nZ721RVOCL7jKuj3nzKzmxJLvFRzcuVYDscNzx5fWwChJx2RvWmXprEVbjDt53+f
9lTgVOrGtJCVgBcXNdRFN3UehDNrhoJoX1uODLsIe627YrhvEai7Xq/ijA4JS6lE0dqE1+tMuUC6
pH95Z4YDjv35MFmjzEYHlth3u84sq0rNHMgUyBJKoszJJwpt7cH4wYpbnWQu37ln+dVFbdibduDi
TJ+vd5hZnz66t9+sIFYjeRv68aI4U2sFlLgRxyH1WwixaHhK9LCFMAq1CERpa4XeM6zNuCWrJk6f
/u6m8eyb51ONUqLcV++bsZaXzucnL/AER3r0hQaXFPDHUJ9+yhPYzHrKEJjGP+2TbqrGvAMp8Zow
3ZL0oaS+HNbAk6ZHM3xE+YrkTEEWi4DDPheBGNW0I2i/aCB5UJu7lg9KT12biMUNgMtCb5l467bL
YbZchYvkXKr37QjOo36+j5j6dh+fQXr7/fqpuFIVkcIpTJPzFnPQAVlU/pflnQfjjCrULIw0Odle
PlI4ojkExDrBgvkP5uxzeT+tZZPqSQnLFE6+o+ir8HcdC5IgpDYRnuJJ+QSockW+X/iCoQS8I5ae
Ud14zkymrWso2GsNutTJdT7/nd81+afLnPftmGtHfTjArn+KEeF6Bw3SWlDU2qWRV4W/hyP/7L3K
nxi8OK/09+BWJTZ0hMdrACS5k9WToZTgGp8JQC0VLZfuQvmboCySajr+6u6WIDZiun85jK/rlX6n
Zky5nX1fp1SbNTuwGo/lt+8tTQOA8WGNmEi47TXPDnJsdPobWGDA/gZXgunLGUDzEGV6iv1F/H2/
dXr0Qyw5uDl56yuEYvdc0+ba8nQlJu9hk2YKR/USQu6F5B1Ldi02FE8AuZ62TH/sicVNIIltCnIE
3knPfIpsGvs2Td5/H9xSW/Ce9l0mYVH4DNrhajXQQCzWTN2dqTrRjKWVxDM7RHoi9g5xzR+FxNMT
RFTGeQQRXQxe4a+1KFbEF8JrKe2AZFSrnm0If/nLzgmtw+RuoRvlQXdO6CXB0tpMj66c0QswoUjJ
tk9LmVdq/MSUi+NawcRpkC7wFCfa2T+hqNlEJ2ZhYwFLEg3Qobk+rozoDRIx916cbb6aXPloilKv
55zLOansbJ/9TUoBCvjmOIa2kJAwj6YE8fjWsZcZYHpm43t9OAysDDEAbe+bi9dQ8JrwzoTKIjuY
9yC7uNn5iEf94kZORuR1b8KLeY6tr9qdwIsNFs2XlBygPf7ARukJsjoH/CpYxmmHwcMu5fL4G5fZ
k14dJPPJvTTGjAq8xgPbY8ntiryFza/0WbtPxc1vqkphfov8060Sz+5CEh82crCcuJ3TqeSQqxDb
Q+MoLH2ooZ2W9SkGBU2Nw0t4YobEGVXqWkQap78DMWvz1VdxthTpByvZQ+exyEIQqRCclehOkPAO
obUM94ex0SWP2XUcRXHfrJ4zluAlVOa9JMyfTjuNr28h3qOhXMIzBz2rExdpLo15y8l2rqMV57AO
x6sGIng9LNaSicdg9PMOMYn/1eh6zRfwkjSJ2TC8ZoiuIVbQC9b3XP+oeMjA2gdewOCJGLNW0YBX
56XeNjuaZYK7x6CZrKn9VudHNYJVlPL3HMPu0uTHjfNAWYg0H4rYCzh435fe0+W9Taof7anT/rVA
YPwXHvBlHhe3UFodKp9erH4RksLKDVMgn5VC6A03D5MB56OdUxtOMRzS40OJjX2BxnXNQJPF8zQN
aKXhJ6fPDhyyMX2sGHrUWhvBDeZmniirx7+45kEwEKBTs0xZdD+0OZFsCEXP3o+yeY/BUkiJnuyg
O4FkhyJyyHl2RVnrw9YICY0lsJVjkKG10MBKTbK4AfEYoJvn1axzZabuDiBVBmjVMAheh3MrtNP2
jmDVG75o1kQHVzGPIGLzREN8i4KU3ONYB5dCtfWZcoi/m9nkFCyU7YQUwQ88FbNC1JZHpmwcw53l
tqY4Xcxhg11HoS0kqL9HNmQk2e0f8VGk4JivCRt1Q4JWEfIZ17lv672OtbhUdMM36VBQm9A0Eki7
3PcPsk40Kbu9A8ez5YszAigibhG2aY6oDq19ZcH663tWdKZ1C6bF9MEWYM5HmR1GMmYh+ifolUH0
GVtH/cRwf6DexYfRoqGWZlzKFZCSdjNh93hf7hvI+QzIhnziODmMGQly9+1aKSXOxYqigedu9CMV
DfkHHMKrHa6veJ7KXgFm5tuqh0T57HefbfPB26C3SLN5JTjQ0wZzhD5xXUMNi+TuPYMB7jEdHDO+
q1LPY/8rXL6whzsoSt2QkPjJ1cXsasUiY2+S0s3+yp9oWZY/aiaCG5OeY3v2dVJszueHwgC23mRU
Pq4JSwoiXFXE+s4sfJXuIv8sRWjlST6s4c/EL+Pn+f9LozClebWoKdhNcaQYSSgWEwY9yy2bs5Pa
UMFMOOZHdN0kCb0nrZkpJe1eeEAo7Nd0xw88JWVzTxu8PzDiLP1rGmJLtG3vxYsiyibKtNH71ZCt
+JUPsfYgP9dhJIOWJkv6JTa7t0aejYONFfLZ14ygb9KLjfvV95riYylJwhsSAHNCpx0zamFk38Jo
DfTmwCf0FVBKmQIHeNARm+3yVQYN/96hx9DwRyM5kISFVUkLaDTOedV933bLhUlrCw1XUMdrnedQ
IriXRsP5AYiRQzCdax4nVox6N2/V7jV18CBxV6Nea7MvjRNoSlEC26qRDypPg2adGv0DgtyZtCAz
1y+Gh0HPAEuuO/q5uD7DXXGdqLIAksw3lAWzbQ3zq0zjRpCIEBKYOcAUGy2DDWBRu7fK4aEuA4Ja
7i7p3bG95ebNWfMjogN1jt1UUd24YTVrAy17LoLk3U3JRd1j0OWtD1fppx7qivfIA3FCU4DK2vMC
Ycml5h1UZJVkPufio9EiwX5rs5jQMWwV/6eOtvn/nlKtTxsDl+wf7Pc/oWO8SUnYUxdlMu4z7rW3
BaZTyE5m6qqNhSOSmLqUqQe2rLCi2k1ly6wPjWgxWhErYVDxoZCsPTls7/0em74fnNriXfPc80eO
IpHtSNpNau6vha5QNKG5JEYMHlhJVrV4NDjxLFHF/v/gxQb7t1sZjhDioYsO6rY0ddR35dyJrWh3
KJJQpnjAwvKyZbgCp8e7cLkaCHVlpX2ezAtxEPX1ftzQvsOsx/iWMlvZ+QFiLJFguv1H+tLCe48P
dxoyqYW84jnWwQP2ld4rjccYggYBXQ6WGaGhTywn565mUK2JZMTeoXI5gtyOseovPKUhhr4hF9+Z
GpnvchySJJlBWX2K0kd0vGMhkfcbGaabCEGi5gs7Qe1j++1mdiaOZMvGXs2T9gaa4C9WVdRasHb4
5yX7SJff6Hrn0Rcb8rhOCmFLbunB8HJvv/cmIsmuWX1Yvc20cDOaCuhPv+ghvM5YrBYjUI+hXt7Q
V1R30DRTun8UDeFW6wiArFGqkUj1BcQhQ55xaSUl4OAfG+5bazuJ8D7Q7w0RUq2x/gOCUpct30+8
v8JJyuz7ESkjQMMQvzAh29Kdo1p21a729kv0iIvG6rOGoIBewuqKxWVt9CdbwmwewYEkBFlODo/2
f5wnqrP+33G7C8dLhB/ZsXp0H8dHEyTYosm91PnDApUHYMUkXgTg0ei3897NWknVAkkypJGZANX3
JG0GLVPCcmUPc0PBxj9WpqcAguCo9BuSe9yjcjBCELoYtQ2xe7GP2YfUAAcKNaRXlEgxo3BKnLFd
NgctekxWg7HgIeDQIM3ZDK9mxX54QtCQdv8xpIlOtZCmPewAH9BLW398jsd/lO2GTRazPmxixgqH
95VkCXOn9BDOBHaytL8MPxd+FgimTtuNjWHg1NLJXthk5jbiOCVo80dURT1Uy+XpbevFhbJuV6mz
Abcl7lxdf8v5nnF8n1K05Yihryq5HH7h75Kjss7txnPmK/ao0rTAohKdxdU+CujNkrg0vMmcX2vL
UiPDXbm9Lri2FeYLaaWgfJickyh4zCahbo3R55/DfzDNQCOf1xPhX01sVHwzph7as0T7CGeNZAsl
w2aGEYEXMvyacCcQaFrTCsjYErpJk8QUQy/hcjSmK5EHY95OGlWbtDpq6Cda+vzUEPW90GyHM0EP
UOQRM5naD/AGwC0sf2q2niPq0381j1gmjNsGzBTlmZiFDJcg7YmuB4rHLsEy24Vq7T4QqHySbiAU
yT5PGsJTPgXEuQCQYAMftFsde1BlhCaKZFJfi5uRnVUZaxkU8yWygPQHQGPi719oTa4keoVM3z0I
3dmmT13SuJxcw15PXKusZKiSot3IUxGkvkhNYhiqcaUcxZiwlDUi3B2OdkMHfM4bi70PUQTGGaD/
pRj5xkUAJs1YAIKUi7M+EvrAs8Fzqlw2y2v/s91I1LCXExLSOgrfDNcUXS3gUey5TXRu2X4Po3BO
NjqpvpiYLw/L+ecHpo4K8bC4+STtgzuQ5NC63SCYKZ3MA5tudTC8XaK3x9sWcQ//fUPLW7mKr8i3
zZ5FzY8f8W7MZpKVzKyNI0ZDthU2QEfgU8timmQj67j2YVc1d8LRVLsHFbjl1phMItsZQ5FW8zlO
YQWOccCCskgp+ANxix/LjikLCE7qnWDLvABHihE/e+e2pakGnB4k/WEK8xW3wEiDN+NXy2ishtDq
hu6D2HJaFVO9VazMOUGsxgk+Wy1nyPjPsx7i17Xjkf7TyKjxr/seMs+zq2F6Brg5dpHNDxuje37C
JH8O0QeAPZBBWGKU8N2Xd9RSts7+WymsYGC4iIlpXgC6v+eo6pWmEsqJoDZrs3KhTJFv5VSwl6j6
BFuD2JEWKY3DjE8WMWd5TYgDkTs14stU3HIcdECPR+OggY7kRuShO2dbkEJWbOCtYH1K1aZhNNDj
oIjFiT4WbTCoN3s4YHt28AQmZErZXeYQcKrOH/ms+fUKXUVfati2/4KdoMrJTdmQ/o4THqBj8zH1
3/JxmdbbmRtEh3rJfA55XO6EIZrHcYTdDHIv+PS9Nd5Knrsu+drXVWTHgB2gYm2OWIV+fY7dVhL8
PcKBltz0LxdTbYVzUH2QzgmKEv5XTeErBczwEocZnOxIvbhhiZleGvsNmSRLipuohNzC7arjlZ3v
b+xlKFos/kOMstQs88J9enyH01yoElLO4D3QpajGvb7kO/AHLQEokDJEzP7tTBzYSsWYmN3dG8e/
xYsKF43gs7fiar4x4/ZuVq36tlhpLbbkuMJmxVSAueHwb1m8RgI++ablMpQmapVAT7aGTbVsp572
ZEakmuDDfXeCTbyl8d+iTfm/OsPrl3dFqofTmXH0DnYNC8IQMIvF2Ox+K5isu1YBHFZHuzW5KQpk
P4X69xS8CKEFR6JaMpI+nZB9Sc8uXvN0RnWBuCOONa3ArgZIkDT3/pEiXPl2ISJscLuC7ULSHCUz
HSRVbtro/YrYdCgOQ9QQeN3PBxFHg0rbejvasN2IPFd7TIT674w2F/9TSG6CvjZlvSG6XlTbLz4t
FWAktbxmyUiA9RwefTEK3LyooenZIO7pyFMY2gd8LIyhR9v7xLBm6agd6n8nzaVqOfO/GzyhMwZk
A0z8eAEZQHgCOOVR6WfLO/OZrsEkgnbG297/KHrVqE3Ik45fnIugyqFT+0jER90DDlKVB4rlvXNe
/N8LlkPBRAKBIWCLH7npEHvkldvaD6yfDQeS+jpqRFiHJxE/Gz0Pbl8Ids3YWlUhKs6bum1ToBP6
jSVWE8itkHwzsnwxugepUn4UOTY+cfLbu626S7u8hn/GXAHYbqEHZTchMqurK+LPI9mAj4SXuVUk
YI/FC6dcvld2ItY4F69RcsYHKFExW36uT3uMAKewzIg7cW4DbTqVKnsr38aTAfygysrvbAfxdz7N
WGIR1hC50evf4J5X5/DjaZoeBCgsCi6+0rij0bbsYVohsazPDlkuXWZOqFlwokegomEAg1b/r813
VVTlhvqaEN+Ecshnl9SqdFi9mlOEpMNXw2TWBGFWaGSl5tRrAimITXl366T6bX1urJ0lWi4gWLX4
zZrK6fPvqC2Rr7c3rSNdkfKgNoYJhJD0cEhJ9KFAmNq2h9Jl3aEEzDtaBnWsclt5yYf3cVjmTNm8
K96Y4+N3yywCDgz3EyCAqipM8PjVCj1MJQPoUpYReNXbwKt9i8qmQxSG5tuG0wV48U8nPrCfIW5L
avvauLVW7aMfSjz8mmfYvAJWsOkELssOGMoBs1ufC+qiYW9/JbsOAZPcxj0LRQtPk8RMPUAlH1qr
yo+5SiE2M2MRhVCsGzkf9tkohZ0YkpJDaAoVqwtVEcgZRvPqn5eOC8xmIkmTveQOgkcnwbuUjcRO
tSkGmKgiZd0FP9H9DMQemCY90WGBpyDo1Xvg4tUzt5X78OaEDQZil2ZqiGYdV7y7yU/GDIzr7mSM
EoCkfTTeUy28fjixaYoGSOR2a2t6zroO2VJQSOPV+LRk/v9WB5DbzXNdFD3+Vn1T9WN8sXBsMX49
Maqs1glkHxXnlRCi0OtevI4RWnSB5Zz93vJNXPkpYzSMtoHBWWvDHSNWqkucAwj7Z90AAYz0KRag
wyBLpiAp9qC0m9f515svVXYc+KRatbBD2xTUcc+rbG+4mVKV1lKb7oUVzdP1pNPGfPVndCA5+CKv
Dho+TVhMiOz4bJLKRRAlhv8IIArTdM9JknI1DHNtUjFv4JgxB7zXKLW43vq/EhQ9FbEfmnCyV3ub
pIjaEygIg5tLGOaBsbN9HpDkJa4sj4NMu4PbiqRSQMVdntsFXNRrplEuzUJFXEKVXV+V65GXCR/4
nNHtgcXqZREIEyIxnTQusal4RI+qOJMScgU2rshbY7/biOIuDbP1u6+S2rkSWkeJom4DRMRRV1ZR
/BAK9tsdUuXeBsheSyW39qNhmEtROqG9jgmvnkwDu+NNjY0jAtQHbiuIELtdmuoqnT5qGO4kqEF0
5z8kacQWKkWSeE1+DE5dibLAWSxPISfIFkP7nwkK93IbeEvf65mu3vv8OlbsUYwNhZaXL8+uEDAn
6qKJ1r9GeVlbcCxr3L0PiPeRA6D1+cEn58spZ+ZwPI605Eoqeps/SqZwdPa/XQzuFOuyn1lRhPu4
CYnUIowi7NXMr25F+0d9ba9eJva0qUXZ8pC7mFSi5ir5udUrojjfMSd5U0HEvImgmw/l3TyWDwyn
oUEviwhUfY0oDDH0algOIK0+VhBYfkfiCFC6oCHFoj3bgAJw/85BjVZG70cG+8bK4rlx1v58M+TQ
u/WBG0ojo0pTCsELdNgtPF4RyTiLOx/bS37GANGvcXbgxCJUXmlSY2qAg6i+VeGl258pKGOh12yq
EMH6wgzRDxr4ASxifr4JW9igvYaDNvB+yJXEIaxeyBWITJrYI4q25txX9wfZmtqToyvQr4wiMKt/
OigFR08P54LWldKlaX6BVRp21tFsLexA2tKqohjFyqR6v0WfJUSSkb6N11ynENwWYIBJ2/OtzvH0
/Jiu57mxOORPLHXlrvIKBwdsvZntn16fIt/DYFdCRqCXTO2SKY6u3c0hxSinxdrifO/Nr1U7vbq3
qHkTmRLypHKidaGyIERPlAMP8qaXnO5UllPO2206VLqfzszddunOrD/wQVRT8A/VkNnNcgcQbbmR
wo4m3wog/88oW1PH/Ssh+zQ9Ruo2LnB4mxGMp/dRnoORq8499r6hl5tfssJPBtzeIrFJQsTyyv3z
IvfkkSstRGpIF/G+btj/0olGb/KO87Sps71qGOEGYIB4sVnj64ZODPbGQaF5LPVKOgWZyuQh9LdR
Ysbf5eIC5w98jKk51/x34z5OdVRd7mn9Wo0yCMM7AOtujlEKOXBX5H2gKTsF7U0K/6xv9Op6vV8W
xCFS5zJ8tomTe3NCpMF1nO/bpzHejBAzorjD2d0ZH7T4xPzT16mgGaJ4AxLez74exOZGdIdi8StZ
RpROXShDeoYqoh2Nf4t3TjDkvWo1W6ybsH0kzzpwibxzL80WkBOKgIAAgGulww9yvHcuNjUjPDT6
sB85PjVraw4W+aaOKYWgqKlp0Lw2BoVbweNCYb/j16xa0wV+xcbu9qbM/CiaCCWgz66MOuSsrlMT
lr9tjNfY6UQC8lAcroZF3cSFj+I69sJiCcgqsGWDvBYaVtVH7ingcAP5aEnvlwNh27eW3SbhVga8
axz85v6Z57JxwWzXm4KlvwDE2evNdW5NG7j3xWvxuhT8ir9Z0NJcpz2SHUpUzvWODRC89wm9bEzf
QZ3bdu20I/akezBtHxPM+Yeufp5MGvlI2YTooIYhmnXCni6h+tDr3SL0Axy+MBH6hdWeQj6TmXYP
2nTRoyap0gD02/qaNhCgTDnRibnkbnejNQ5KE38NpUTXRUgC8R5iNZ+if1FDNujLa0Bm6zr419BX
F2Lafwhp5EBkf9puw6nKkb1RTz7Ffmuy3/OFKKiA5CxfpSgPib/obUiZGSffhURfRfS71idkYTFQ
znaHzSym6j5NGYCtHTmqZk+13yS67F/6F9GiHMiFFnZuJWO4r1Qs8Zwn0RbzbBXdP9yxAJ1aToFa
Mwh7nUVJrR9tGe3fEJy6IQyWNUE6La+VH/qQMY/wpVLvdwbXx5spQnj+fYCIy/TPDiMrN7wJaRwQ
oRP8WBp26iioWaMEhL8VFS8U+lL8vm20f+85Bb5m2a17AkFaMuI+zt1GkvOyhliAcyfwzZ8xN3nq
EV1wGtA8rAyaSqfkCQeT/BHic16CIwW+l9latfGXpTsMpteokG9v1Plg/9exbwPHBmQMDgTSm+3m
+D5EPkhEaotSO4oyZYHUAb1VgcesRpuI+LWWJuYvbtIPwYbWLj+QYoKD6KF2HO6+tn3dDj5Tp7//
5iu42bjsvf64its2fwA4yY2J38zVcWXAPC4QqgscmaGa1HSb5GQhlhTrVg/KNHoJfKiBFjQIlqZ0
OtEkycXuYOlrdaaa3tQNV/2smrPb2tTFdSLsd/+8MnnPvtUFQiTICagly2FLcolgXDXJvH3tgxkP
OnEyHzvpMY1Vj4WEgryvY0YNR0u+7IbDuzxW9g77q4d7hJfxnB9BjNYZpWC6Z1M1ksSw+Pw0mKEU
G6BcACf1m/KxzQQpys5Omnrh3trm8QJiDzlDIwADlojZb/boS4KZbnfl131uhGmE7ehBeF8tpUax
NMcX4iRsMeJnvPksaNXAOKSbW/7JL6lBThsLXvg5juFZVA20JUrUkrei7g3gk/QkbTIFtlXwjLE=
`pragma protect end_protected
