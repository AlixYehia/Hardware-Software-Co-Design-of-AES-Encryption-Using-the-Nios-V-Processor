// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rCqVPI62oI2+PZf/dmeSb38H2H6aQ4lAMR/WYYWL0u1wTAJaqZkjULofYdBjKQhLKT9DD2GgpBcM
DG3UsoZfciM9iycGsQ+QLLuIP9kSfMmzW4YYwfC5FV41SpgLv9Ixc6V+Hf7yOoFA2KN6foivcEqq
6QQ4WKljGp23WKcXotb4FP3eoy0vaklOCIqCn7dcCDbYpDHJxDnIHXcF4QqLS7AjV5rd5NWpVUDV
KqEQpYvICC+AWrFVhDPybpiz8EHqhg36obHOj3L/buYTDD81Uk1jJ8O+w7EeUDLtHJnTTpH//bqM
GTUpQUjVXCEkFGaptujb6HIjg2HVstn2vNCvEw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15888)
hEvJuHzAPZ/V3YjbZBAWDa4O7uQALRzaZkX3Muo7lPLqDr/SZAW8C2njAff9tCyGStFlGs5hKe7f
eyxNrQjdmXjl807g9IcJvFfKD8zotmTXGmKO4cNCo+xWVKmqgpwv8pVqi2fAr0gWzgAX+o8OWetD
PiZggLFYwgFHIJLY+D0ffw6EJ03mB+CDHKM8NYheeVgkN26z42bDcRALX0Qj6wwaLnoP2WXWybvr
MJEafTwMPmQaY6GvDPqqhsVlRZCGh88klMbnhJ+F6LUPoueDq1U5TFjxjKV8WzEIPitWogL6L/rK
+UiEwV0LDwfzd76noRkNpLzbP6S1tMLYwnMIragG3VzKI8r4+VOo4Q9CRfbEC0VCnu/SWo4jpQjd
Fo6u0Ue/M/W9vCcgOMhMeSkBzAnQmpsOwpYbm2bzLeLCEOAb8UO49ZYTEJooemzyNpVGGgpi8q5d
ywzqxzKIbWxr5QOn+s8BZFIALNdCcbcwOiFHFOFnV9fcgYgw/M0ciShpTT/bnQc6CWN3eNF/H0JY
8xEjQt4ROHziMlPdY6YTeWi+mNqRigQvemzblMCRQNc3o8qErSwLjWVRFf9x2W3Pm9ErvLT7jP+4
jtjXH3pawC3IeEcRGjGuiAIRCZ2LXChTs8Ats9bkwECuxDJsNBRb0Xo0YKaRiyzjIch+SQpMKAQ7
3ldhe4tQ7vMaatbx81s7kBs0S45BGQdkKUN8/b3Zei49Qmi1vVjabAV7FZd4A5x+tkBGnnvaBiB1
ANq8ZquzGN7rFdT5UunS4s/yDqA866F9J9+wXPYpL15rOiokahQCfRYWy6xoceo7URkXSee3EilO
WcQvBIo++fJO66W8Kb23ORiVjf++aiPqduJzFjQ4nUdXjs28fiEz2KK6Vs74Jyw/c3uL/hCpehfB
Rcpl8MFFv/kzSoFLLIlk+BzNBsA/d5CaoikuFX4T3FjdwIvJoSDY6W/dXyJBEqgt0jtJ66cQJAqv
eqhPyS4GTDtyYIUb8k6zPQPRFxAzkQ1Se1W2MXPK6BwqmdoiHes+RMenxpnFWbEaMkyACgZdmh8Q
4lxIPbPrQZIv46vwqCIkvJeHqoLBFlJYJnfnKM35ww3LnYlYXoHUVqbSokd7vws3oCqR/5mt03g0
TeUZBbpD8TsTUssfzj58zxB8aQDVar5Y9c1qKSnmPZjgplMFPd8LC4D52ellDWNUAa8ZCLVhY7tW
mMzKRp+NjgcujqfU69xf1x3eOHv7mM8tnSlaw6eFa1tDij1n6dAygX/O/mxR13hNPFFlHcIu+wOL
Dx5FMzWFWOj4s4cC04ThL9mX81g62c9tIWoQx293p5zsty+LQ31P+SccirG9uARuSA00O3bUdpyQ
y1YWkLEj1phCP1b6Lib3IL8boQDXy9i2zrcLtK26fDjp+Xrh3lcg41F+lNycuKp3zf1y+vm62MWc
u4Em2hFnAW+R+rN42t+Fln9jhoM0MXk8jYLhbOSckEjQy7yeFKMRUOnIMnu4XoTpq2Md9s95ybV6
HGt8k32Ix4XxZywKylgqkuQy5GqHqtjIp2y1VqtYt7k3a7UJeZu7t5YUfDerLrXdOiCZD/nDCC8e
ufYiPYTxKiblO3Kj88IBcqJSfUleJcSnQWUNKM0o6X9anf6+FS9cBOundlHxKYqfjjZ/y5Uw93B+
4qVue3MM1QPjE5fL1A+ZIQZVcvSKAAb1vdq05iNm99Y9pt+3grbdVspm5lU4lumFJovNUr83BsRC
VtUzxRKgFbvva0wawMxTneH0KKvtaDdA1lnY+8OLGMr0u2SVrTPjVoya0eLAQ5w4ZnvBX7o7KFzQ
ZKOJJ4ib4IOE65xJryGLM+t66ZzlDZCUrFyaCwQBqP4zOtKf4A/YidJWEHgafy6X5sz2fdWIHq2L
SJeyHMpPDu3fxOl8TBw5UX2Byb2dTPx6yJgLZItTq3B8/1Ln97y1iqqd50lMiI9mkECIAPK4dMva
F3lc+Kx0jWkN+2EeV4+PsQGwqVUYFmILHaIu4rNkjsG7oN1YwHv2IcqEcfa75eDwvyRZ3RpgG6rx
gecHMJarWuQOJO9MbuPTdIaH0YvaCymfC04lyT7iMyyiZUmsrS+v8ASdecXftk6Pm5T00c8uNkDS
C2MvtoBNAaBRUxK+HfspoOtYDDSC+KUUeiR5ivv9mbVlyKLgPCupikJSLoYFYrNnTtN6yr17tMlL
DK+D+wtCCuAQiTcgfP/5iFOK1W61rBf+B4+bmPZMmt6Xze3xHCKljEmCxLKzbY//n2jgCgE9FC1Q
A2JaW4dlQfCD8K2HsunWLyGVH3zWf3X3a9HIBJUsDFmgCm3UH+dy/qpvlqQScEFWnQFg5HaiECHq
RC/ZEkpwcsoxHiIX9Bpve1aphDEgTaGPoQ9df3C3pC55DXJmcCoCGB8Cp3mfxyHIpRaogfYzzNQQ
iYf8V5Ab0uyUET1hF/8X9ujd9ol0BfuxhWW0ngieoNSoIv8DgJkzBF7YdCclg6Bf4/NRsutfAm18
Ps0E/R4FhufaSqnyD1YmvDEs/MotIuwIMlAwToOmBJKqEV1MmKwFxm2CplGoFLTU7ew3hTUn8iyq
SVPWppbliSMldUk0rEsYwEBLXWmcEkEJYsCfdcQt1Xwdz7Ku7WWg7UR2gMHPZ1sASfXuyKRRMLYK
2O6oTwr7+0dX43it87UwUlyqVSstFPdx3MfVBv008pDsALaly595gEdCA507ed+ifpMu0HhL/6S1
BonLQNwvmc47Y9vT9wbV8VbNpuaNbNnB4mnXQRetuPP4o71unu97csJ9PTf11YoQb/MsNgXpHfLD
L0PQANVekS6LVhw5fv+OLkSQEJ3Hi6d+DgNIiwGd9gFefCOr+wZ3yFhaYXoG9P0mD5yKdNoJc0XN
YN0ZCee51UUIM+Oz/rahQULK3J7BgzYYng0Q0JJ60qWxuCc5r8j8z65SWSdDNZsaY91gWyecaOeX
Obq8IksAxdyOeOuuGPwiLgEIjM0aE8mt+g6NN9cClwBdhLsVzEK1yFxp1RfLvC9PGKKpPDvBVJxw
BGNJwDDikcaD8o87arCzHDfHSc1iLdtYJS1fYcJanUYw+HzcF0GGR74sb3f4x1B90FiGLwoFd5Wd
xUEjI5Bw2yVmPvX/VCqtEHAFjO+3FkTFWxtT9Bg+WQJGAdz751qNBxzngu1RXqQi6NvA2/CiRZHr
oyQZtqEMaxILC7xXTFXir9hWckc7gEZ53Ha96+t3tnMscfOghmsXUvWrV3zeJS3UeZJq3qVKbmVI
rrw6iod7GNhn/79iHhXGAKuZr/svggcscN/r4TyNO9W/X9gramdeDBjFjtSTUuKfxQgKrEbUd7fv
dtPZPxKDnppNduRkdBi4l/UFaOR/HbJ2/BQKcAmV7qQCxEYvc3V/YQ7OtTq4yNV1MiJPwffP+NuY
31ZHR2Kq5Rh+m94/oXI8R1OvkSBtR7gFNU/YGMx3X1YR71SmTJ+ym+/n9XZHh2R+IoYF0xvYTlNA
i2CxcWk2iEcf3k6oVpfVjye4Nacuh/A30SXQ/bFybTWaRDh9NsGBOyZ27Q1Sa4UsjwgJTQM7nkfU
y1pVeTJ5myd36L/RP8HPsjyqX/i3TPy2AxafwsQIzbbTGNgS8CGZMjdgQXMJ0oQfSWMSV995N128
QHBi908s/TpgSS36BU6T8uouo1A0zIFN/U40tgLpOcSaMn9CqRgB5oL6XP35Gs09F0aXGn4WUoFM
arOLbYgadPQb0xOwi5gcGW4lgZNgCpRlZWuRpVVNXNXp+wXU+fHzC3l1aPGSR763rtxPse5BLI7h
tqNqlHE8L1lp0VD9W5gWmUyJYMA2+uaC3p1O6FlYfy64l5OrdAhvZrEP/onDWsc6hhL/kcQQogj8
81qt5gUryC/VwsXHN0Hl+EeKXO9kYQb2870qcpjeMHmPtfqX9Sk+H4cOaAZJcDjLFooWbmjA3x8Z
anAst7IsW1j9khtuTaxCi57dYgo3fb0NgHRFhu8NdyAXxFNcOERSpJ+rnAB2S/N0lJc9CdtsARl1
vY9xfK/XAlUTU+bIb2wBgJ8jyW8t++cTjhTXbyaFmGGCkms0P32BhwUlmAxmBAP/E1hFaYCd2Wn5
a0nR6rVcFgHDZjRZTRsLjMAx0v5XJ5d6X7DyLxi55J4Nr6WnT/qM1xYOeBSXbanVNZsSetQ5HkES
ikt25V7deYczPYLfSYL/wFFUvRnIdHiDCeNObCGhP0FS6FARAsWUz50lNxzvQ2Ao3Av6g8gzeWdx
QAhoRioBdcSVp9y1+kRJlFyqqTKCNqeT1pRR00tWf/FGcCREPRWrE5By1F2bcQLFSxkMI9wQMFLu
5l0JESeuBBBPvZSFEHFtwA8KusaJGw70YrViIGqyTE2vmD4Z7XpSoDeSzma+5Z5BATXTBtnyA3oc
8QxO9vKC2LMwKsFBVYbcDITjC2mMQ/6fvDzRdUGrz5mf3vZxBRDpeU9tO3t5zniZA3+5un0uakKU
UUfJf2mylc2dvVm3e9TV+iYmCWFApjL7ittc4Ywokkao8NepbAwVD9JfguvLVIYk45NDAy2fIyez
CgB2FkS9jmRDlWnzuh+dMeosD615D8DXW247INyWbBxqFONuAUsfPB8EkF1pKvBwN0d2xp2hgD5P
XbjEPeyffnZ0MV9T3KvPIvvOvMjmVveYUow6dtvLKXK/Vh4ywY7Dbhjrr4Hs2Qz5rZYgMhcM0YPn
hCqIHgWYfbSPdlr/+l6ap4EivW400KQnF7uXTz9bPCOoSMaE7PX+TifickdJ4fbqnlOxgwCj1ym/
ae/eP3Ggu4g3zsIUYCxXbIVL/xEb6+vwfV/o7uYa78H8F6j7OIpuQalfGzwmtz1rGMj0m/IQkzOK
WATSB01gUCZc/yS52aWbviq/Oy4atcQ9q5TjAe8Q5eoU2WXPkAFFLqhRsoOMD/Wb/q5o/Tl4agzu
RsBjGBU4JUOuynPfAHXGHTjTzMgC4hCCvzENsr5VYUi36LMl/iyrBDJw9NjrKQ0uGjS9A0S4g94g
yeOsAJ9pcwWxwuaVQs8NggjvOI/kpKNfHxQumu1BYKuTsgsk0/KEdBVc5MK1shAkD+u0MrmNUAKH
KqlBFY3qiAAM/SuSyjy6kTRlrqOM9J3kJu1zUf0uNLTBmeDAxcZLda+EOrovmvnrAvpXjET5mu5f
Xg+aknNNAKLodHD6d8voD8KsImJiUNhKQnb8GNt+U3flGm5tFPtsZBDAzZx9DlDAk1u9deIV0PB9
hTLqeQd6aJGkP23uPPATmZsUJVYsSmuDkaoT0VZMVoPa314COYxmmRgyfm8z18/bWCOHngdwdi9Q
fsJk6dma8bKMKcC5xNfind0AGRZdkr10ud0jh0kIa/AyisYrbx29xtsg54CSvOhKzqxe6L19xjbQ
TyQd+wZ41Ir75RRtBImu+RsV6v6S3B2hE7un08QFJoUYdlclN9gaMmVdYVuGSLl+0xK4gv0LxY5w
XaIhW6BXrAUeQEYrLZ2UAux4ZftLJ7fTl/LYGMJexshj61+nZiuHNyami1GsFNuWdmIsHjA3TNTG
3iO2m5QZGylLvEXjfqwLsZH1OIRWPNqUTEWqQMvUrvl+DVFDioeCK3Q4dMpMq6hv1aOdoVacR0Pw
u8cZvchE0gE3KDHfQ0xcKmIUv1s10iR2sVN8VJ57rOn2iZscBPqe1SUtCfe4cuI0at+BUw4pvtB+
FMfQBe1sE7bGHDD8A/Rphv/Me4mM9p6xz/tMHWzie5sWGN33R2LREPFGQ8Be8m+VEqpsCP/2ZDbL
r9Hpt0gWngfs9Z7/v54XqF7MFr/okXOnpPxWC1bGByh+PViJA8PERMt5KqXjb0Zhn6Ql+vNcvI6m
KAQ8ju+saLmGCrTfuCbtDzsuPY2daL5VvdJN6OHHBxSvIkvHoHxRP82XTDmqBsrsOO+V0k1AAq4i
1gnFlAjPeNHgebrTTkSpB7UmI226V4SwPO/YW6vICYLozI1lf//Tazs4zhNkmyx7nF1mtJ/KglMC
FKnC2qAMdJ+7kHsHqVhYbDcmuaAb+lfnw5VVpceiZWJUtDKRrOu/TB/gXhHMnvMMzPN4cz7EdcSA
vKRSdAc2r0u9X2pefHx1eDdY6M75uHO9KIFZmWnWp1T/3Rxpe8QCT3XwfwjiAtm2hezYvHoDzKFf
Xn/rOo0/lkGCpkFyF3GXrh73QsvM7KNcT4genXRU0zFZ0tWImhxBd3jbILCplm9jS0OgP7ofM3Cr
IFgvUkz1wCInj1j20BZQQej/FnP6+o5wVBd4Vo0IGR8rtRM/4hncHHVHXFIshKvVJerrXwR5+RyE
nmvwENA9FVtsrlqJlSsm3SMzmPbjhQkQA6wIqLY9LY1GGntIjgaFRV0JehxrcZGEaJiaH0sQoRb+
slmKeBZeYMsFB318BS8w/ruVTTTuoimg2Tmlij0Hzp9jvaQ/PEk2f04OwOBkLxlxe4wPQgO7QUmi
ep6+FmfsVNKTw4ljTJcs89wPB+1heQ6SsMr7SD9Hp8Bp7OfocGMvLNXI2S7iE7B0RMYKVLvM4+8I
uKwBpcT7kZ6pQXYhOHZ7q7dz7tABAeMY6UavFSkv5GkakL+PdOaMaysFX+UZtgtPpEr9ybb28PbC
VSKZlweZ4+noh20va7e/7NWAPesy2RTeSuGxkGNJg+FdDeBkwJxvnE36OIctz2ZEHIOZEagjcI2b
NCX9tEpOHh0nTVYsj3QbzXmmjBXLwCbtrC7Y1kvDlUzWnkZ1oKQqrnQgeo0hfav/wZXlniWFzgk4
ZEIC9JT8CxPZXZiL1dXEgOhagHp47ppjVbNZHMdWBLli6gyBAxPcIVJeWzzx+qRjNoHUsXZuEEUQ
6Uixl29cLwSTRetxQ/5c+W7R4CVyQCPbXvRWE6TqU5mzcZSSOxL8MJuEfynqy+yC3myCNCIF1sfM
8QqROYju/KbyrUAFjCpetkL00vhj+ysqnH5st4cl/9TWvt5N3i6zRowuDEbpsyKlQHGrnBIiHxfG
qIKdRRt/vQ4HyFIYD0KQk3I0pBraXkTvh1cARhZdSvaV8qKZNUZWkOJVeQkai01sWB8BzTNJEdF4
Xlgt+4GC4J+4icSFWq2GQ67WjvOu5ZWvOBGM3xWiFhQfwP3fC0DPknps5Eyp7XybqXKD3n1qcSG4
8zX7D+U7VuwNgQGJPxQftvixvxlEF40zphjaVs8sehESzHzj8U+jY1gw4ZRimQMeeEmIr7K5qhJP
ek+Za6uhtz9RHq+LuejAnRZUeSRfqyy8h25rqSeMWZ7TuvjHRFJ1Af3obaAuyrntdp3yMzKLEbqH
yNCG+H0dWSTD+E+d9MFoWaIlyqbDnjhUcqq9m7vcsbHUMQ3VaVf9gJpr6rHOzTAW31+AE9LDW1bS
sCKpuExe7HNSRZ9HBBM68ZsfGFfV0ut/wQcntpaSnSzKTCalqyjoQ0l/UG5xjrcfa3SaORAQft3S
RwzL76YOYg8EAtrjXM3znPXz7CAAAMSphP3+Icz434AU/ySF/gZrzXpsD6d5WK1XgkP1C08fLZxb
0//5GWNPYsQifqQSLXEIJKQxkQ8VPyVh7+7Dg5yU2OH3BisPI7sDQXbkO/oM3Fss0n8ihz03Z5uq
mA7qjI9OE2av1UCeiZSmLYTmyq24hWqqoqolOqy3JTYw7XzX+Mjrrtg5GnHrlA+eQkwBnrmE7rOb
hvuzFJwKieGhGxf6MYxzKhMtL9jBOAnFZ1if3rzZa8zzmfm1jqGajGYrIVYSs4DdiOpX4J3X1L9b
1m0ztew6GIkKq0v5hQs5Krowd4goZ513SML45yaF/1/jmvDdOiXlnhbFxJTYDogxkxeyHO2RoBZo
EjtAEV9pCeSJcZpoK5ZBOK1Mwy3tDPBaUaUGV4CHEsKrpX+l1MsEmku57u1l2pqoIeOwRPQIAZTx
DQuumOYC+LgEogYY3meLLmJI6/ISDeSd8YX2sCl+tvWWYQf3Ju6gKPmnzQOOITWiAqjHwWHuVwp+
gICtqWiDZndNYk1+mu5mflz/tnbxTm88QAxS/NtXH9yPB8zFiahwXFIUZTAUx/EI2Z2ULZiJOx0O
dcD4N0TMrW8qH8gpGwOy/rLv+Ia5dAqhZshFyJenyOrXY+fHO6TgHUR1pjWt/lzsx06fXIgdCKbC
XtUm4OEk7GhBTyqJfJ0z53tugR9Le/42GVPGkFed07+sqfan82r9j9PCDyc3a123ZcKZkjnv74+1
W4qJKwfJiXtXnnYf1cLWFqkEj15RpmQy1jZ+/XVdqLKoCW5iLC8I98zUwZWZaLRV3IhWlFm0ePI0
Jf5F5NQjsZWsARw6fjMDKELyDvWLADE4SStRrZtsFRuhBrM335ggdk/L+6CbDByo+cAufBnJWmXA
Q1+JXC8+4vJzZWQFw63m35I98P+x5WUylfzgWivK89mEXWuJ30MmA1/V72UDA2uvzXMoXvxn2RrK
vKfXlsssYefvTzDfo/NM5BipF1IsZYrQkiuNDP/Vzk1A4uuqOgge9nuWA4BBtikeNF05jlJcppBP
hUNpMJmqi13KPTQBhQXfPQjHtkj9J+XYdNxvtLMt/nRBafmsGZzEV8zwmkn47JdapN7vbRi3LB8H
G/B6ZkTfxHk6i6vHuF0qSZ1XyUynK4ChWWHxqJgcwIDvpX1l/fzWzu4ZiYNngopWWONjlJ7ct8x0
KaBNvcCqBeYBpfgVw/WgEfRnE1m29Qk/Ybyfa1vBNASyWvOGdmgvvMnH0ASHqCSEngaVDr7WvIXx
0eK3GQwFhKfKOsGQnKXdF6STcJRTFDDT3mgOWe+uuVL3R6xjktwn+UpmXPbLmxr87f6PHzU0QiUt
wvdOv3zzDdjOwxhbu1wXmVJQjX4KHQ4qXo7z9EspNC4tpaOYicseFH6j4W+6OLV38TmfeU+3Xpsd
3qGYDbF3O1cSJgw0VnRbsRKxehe+/pgV/4Vs1qV1JeQOcJkhDLXFjnsJnThxFNB9igx+txRnnpdG
JdyYem8L8SUIjOrycn+iuBM3D2TLyYR8nvG039vqyChwmlcELDaMaHCTTf7b9FqTpbZ9JSuyQWX4
Lpq/osxULStbamPHG0S3lAuFsOyPlS/nGQmdvc45sbzD8wg2TtOXtbV3honHFFse49xpSMVUCRt3
G+puV5IWafFITR/lDCwBvD25w2uuBlvVBCRkwQHBxMkVT19/QEQ2+2oD5FJVtnorKq6iYUwNkiFq
fGKGG3JxJ+2FDt9+pBxUgMFV5IwiKvk9f6A3ToZ7kcfGAZC4QDDZHXnc37qVtJ02ud+FxHJhU+cT
m53NZDzA7P25Xhr4hcb9mxJSgTNnwTPO1eRVGngEqBtX7RlG1yaw0nxLafmc+y1OiQg15dws3Xan
g8NjKYDkKQkCr9ZZ+9RD1NvwBTMQxYg0sVwW9iw5wWmfmAN2IxVcmKqQ/5WhjFtQeb3ic+6WXjiU
2p38pEvkqX/Ke3TGnU3fBujvuuQgpZK0EH3u62Z/YdE4byb4t/F+3AmMuGye3fdYKB8qtReTQRis
RaOkdqcEenBdldpjyrXJKCIetT6274XZx9/wXWRHCY0mETkPpWKrOTpHHuwM0/xyJx/0QVztU/VH
XfpfINfPA967kWIlUvBHcS/8w+z63h5iB+9kyU/LNZIRunvM3QW3oR8AsGrOVqFWCMSz3UDUnYd9
ZxQrEknqQ+4c/kOMQ2XAp9WmaCXHjeC2f7GGdRPbeKOf7h1xXU7V9GnrBpnBuNoaZPPIcw/qUQ8V
kQt5Yjti2YIbfn+cWj2mFpKKV4Ti82gutUIrptVxjNKHTCVh+lkl8XI7a3QgmKmkztoS8fpWjcfU
kWzsvV0hQcPTKFLk/ICUaUS+xJokYzruklgXVU6XRAFA6Nr7E1hcjWaBSE0mD0A3lS7GfIDXuVa8
Vt8mmcuoE+VseOoDeOW91o10VPkSS2UieUK7etchyPZ9yhop5Wxt+LWVLYAFmodWqe57nchKGVNd
r7br2etC1flj0X6lMM+xelrCQSXY4UjB+dxffNQlqW4oYEIxWUZWgrPWFhhvEUH7YsAR8TOGVT3r
gZp/pO0eaYB3gfpTh4wqb4T9LxjZa4xzlMtG7swbHgAYKyO7QafPeNv6EovLZAOERKerL6XlS2zO
DXOTXHoCkK2+SEeyAdj8UPkq9puSfhWAbyZihGKxv1qRlqt7pD1HPLgg32BWsl9HTk2rtO9SpIyq
/GEKSaMnS+cPTIz619r60+UfeyN4I2Z8Edf+z3qWrtpEf2aKsZKz031XlpzS2V52MqWoD8UBJYbb
OqJYwreKQzLELDKCHYzDa1VBCfMUV8wqXynXU5L1MsHC/Xl0SiL7x6ORAF9A2OA7Ek6taoqLVnJM
0R2CC/uNP35QMQDnR0kHjPqKHsd6Wm3BEK5yfu+OaK6UCMiP+Mbc/PVVqtPh9LOwRB++7y9hfhOE
q3jW7f5xjOCuaTM6Xz/EmyPUrPO4fMIxOAGVI6mFyEP9W5mRYPahDaWTiZZr15By70unELHS6a2W
Us+A+8JtdSMvFk0XzzPgDSRhOXWTo6ahXBmQb9TO/Ir3pSKWGDBdPbaX5ib4HFgyrzv1xHJnI+R7
1q5KF7QH0a0JmIVyaibZjOhBQSCoMKerOIgJDXTWlayioirVgstYFUtUdqVKRJDRC2HWw9SzkE7E
NSeJMtaMsAlPy7LE9cI1U0f7xpcnyZOw35eOMniC3TTE1x4kz4tGnYO/qojoLzEjgUGYhGujpTif
1pJp/67c5mfOsWifCKaFZG389qy1jiIlpQyTqI/nAo4+qRbZ7lRWfRwfZtU7fm/qyMInV/Hv+ZrK
3NkI2TWkmlXgoRYsQteXOeQeHRQKfY6jTxFmmb4Ve/yeBdju1zDPJckYXOTQLuF3+UjQWCjYbLfN
UuHlnFl59GrgFmC/Rioyja+GqNFHRA2IrQFwy+hg+cuZiLxBw6OidZpd+Gi2a2K91CvUfYL0RhdG
ypBLbaWhnZpOPX+vpnkXzOh5pRmA8Yyw5BI7HQVNRrKdZNlKx8cIY9c6jJKbmOIKmuWnh9hcOPri
Mq5tKh00+m8YqsdULdKcyM8/ICGl35VXdCF3iYBbVqDC84JBbNhXJ3UuqX/HRazlXvFXsIVenKH1
viR7ugzShNDS990vBMJQQTl9sC2Q2FKIeyE7yZBei+0aOhbEXK7MSneV5qpFWcOM/Qi3Wx3cebvn
y57fBXdv9Vsgo4CoiCXh9LMakQDsuAbnqd6JG5sycYiRmQ5aqetUzw3PpujymA4HKm1VuZG2PQXI
6kDUmMpdBHbtLQzrOwWLCTp397zM03ahyYpesJrTLgUr6XTgv2M3HuDif4uJrDgXhSSJ+JMH+XfO
6PUSQehY7RkLNAhFu9GDlqfcCM0dHigQHESQDc9iAP6uuKq8Z/HxrQeB6rU0yESkiLDncRwScp+h
Jylf8Jr+zkPTtWK1/jcBk8Us7yUu+7LC/o1fq0cJU5A3pbCxLZq/dpWXDW+SR3CQPaAwMaCq1I5Z
VWEkGh0gAty1gZmIsiGka1hIkc+2e1hVb6avyfnrOnIQ3tWQr3Ee1vU0xRok1HlTLgo4bzOKI03r
x8uKg7DIIkS59Fj7RItddMtzENNXCj4u6BMwrMjA+BYfwssRs1OJL4QBExYIraC9/YMPsHHbTWrp
KLemgrljqJjjWrMvcgxz0kGlkwZYnKnlEKJv/KD7sKIVwBZI2QSrtXUkJT/oDExHr3FrnTSqFc78
yqyscFxQo3qijzRzulAnF6EkHZsNCm7agkA42PIdh6ny9yo4bP3c1Bf2SPLvsHYARyMxWDB8EiYR
XmdrKdqA1EIRNsV2xa9F8oUL7b/akMghkyZy7Egn4XxdhiW3/r3kFwJcfzI73hbim/lNAvh1FxVf
jhKuP/IxTdMo63LFRs3Hp/YR62nA/o2aSvrYJZvdNEGNj7ciuRQ/pPiRZrA2ELKIlCeNaW6EDWya
R/lOUnOo+k/s0wUHxlf2Z/HlXiy+19ITzp+BNd2hXqa8zTq3RX+cWSZsyjq3A+pYicFRwIqf18C4
YTZyEidF0w3VglVuZjYPnXMqTh2DjIs63y8Tnx87bsNGOkVLnfnEcG/fFWEpF4cDoT+D6tqOv654
s+mAwiwG5wHeum9xvTP55/S/LQ6+ILpm4JBH5T4b569BrNLf9873pnOyRV8oBgI3JOTAbb0Pwvba
rqpA/e4Z50Eo4CaP96qxtK48JgNCimSnHliv0IweCioM4/iMlpPvLkIDl86r4OM5NF07SDlPQ0M5
9R321mNZg3YfXM4fx7utFarxKlZG58lO8G7Sgu8mazkgttzyeLYhD/m6Y7uGw0LzeKILeyJtMcbx
+jtmgn5GrNhppqAMrXcPbZljYlf8adxIN8esKKkNzxUy66G4rPXLCAzX4KXv+fIMu5vIc+x38PX8
6ReZG3dPc5GssW5PjhxLr19Xr2Qm3SiG51/7O0LEvnayVGiPGVRbh9Fc1F37JQc/LYZZFEnPW4iF
4GA2IgrqoyN7h/UEutxLWAqopdbSQlXpipc8TOnttdwmYnGnBkWdKfaVQo6768dr0L+JErSMT9sG
tEdmanPVL2PRerafDCTOr/hT3XcIxPuzzTr18gXo02ib9eNw3yH6KjM72vJKkqV0xDgwLEtfk48G
DfGuAe++Rl4V9Q9L6pdPvs9669IWFDFN54kevNBY6xuHis178Q2fUQY1kHWF3bYl1vhNTZMwrQ0V
DmtvesR12pLqbkuWDi9SzQY2JvhQJ54eIxY2/HWx8TB7zxJUzh9EfhbFMV67mVjk2EPsob28VjOE
ia4K0U+0fVyG9ajC0UP79JoSKS+x04ZrbwTtWVx2HaPrG0OHG1aK74Yv4yZjRFZ1K2PJ/eLxCneR
hhh9WrzJ3yr/zoMIYGvtyJNDvIl6gE98JbJ1TbkbzOt9/KRh/J91DgGXEgD1R6hNghyUQkNAZeQD
xiFHMgxNjkLV0pI6SbnhZVaVIgsCB39MehI8fxjhSBO/EeIb2ZMuUh6EYl8iIu4uDH8dYcfWEDI6
5vmoR/fvVkwaGq8DCVbCbds8yDjbEcveLuuoeOi4MlS8QNMVS2DGA5xJPd2jZdLyq7LQDHd98tch
coWAH5zW2JnJd0v3b6GKBo8NUo70Yz4gaJ4h8P1lv6VWLhjT6gt9ZXAfkg5S73GzI+c5BlBstRg0
UJe2jRmgAd7zL2pX+8cmNdBzpwaHgCQIQUthEwJk5DlsDgUepw88BdbK4/kFwdKpFWWGZqxKeQCV
0Zh1IU0nS+lYYz8GtFHpC/+CiI8Q+e6lKCdkSUilSHVrHn4yLqWXDGNIuejSMl6ZEPk5nHhcLMux
xMIGNhEdB5zhaerF48DY7XafDDGQyjMmJjkZfQn7obKSDM+wZGMkP3p6Tzyts51TAZ+w/plLwhPa
cMxfcMtqOEvzYr50PPX8j2XrKQm2/rWGjDMnLjLbw/3C/WziuseHGvNCLNQJbXNq3HXYUqw2NPiK
0lhnRO/ApyNQ/INYg78yx8WxveSLo0KIgeQu4ScGYay4urig9qtlle4al9qPuDD+M+kMOZiVm0NX
jwT0X3RQhCsXG8UnXh3q60r3skPlxrKVb301Zq7Qb3GoQfEmnQI6MpPJxARvwVlQVOxKtvko4LfZ
VsakoocJGcZxQ7KtomUNCHKka/WRt6WJtQFc8StWJUHq0iW0ceaV5kQHbF7q4ALiwjtcKmiPRo+z
xSNsbXc0lHf2QYSYtZ+WMGpDr99yR/v4wPjl364b0WbAnH7jcOQdPKGJsuAjoAnFCCvcztmKiUpu
Z9Ic5iccefgGYI90AFtqcSQwuSTFDCh1wwEP2IziGxryqLbvAW8bQuE9vm/txyBNAqh8jvf8dtQb
X4sqDYgCkuYaJPd2Z8Zz6klTqKoN7LT+0xQYrYBuHuiMv7jMe/lV97/Ybci/WKFIKo0aFaLZodMr
cz8AE8lEFCJHZc/+UdXjTZSQDNBMO7ZygxgraZWotdABoUSTj7choVTiUCP+wu5sLfX9GJtkUDx6
Ksma9/U1JWhEdjXB5NVXBU6S/kcLpNor7VLEKmINZ+0fUVVUBoFlXmyx53R6A/aDH8+NhpGdmODG
kZRrfpA/2uPgNPjr+dvC4lRLKb1Hi1I2JYBvhXJWj7O1Nk7tZilURxBT4NngAbc3UOgjbjDkrRaS
siaKtNVaamU8bJJ0b/flnTHdWkHdwMJZTOzhD2PoYufDjKdEgbygYisnHa3N5J973uBJc4syciCc
vQ5KXrfq3XK3tkQbzCyI6wzQjk+mFv1PAneaWV2Cvg/mLOcPxa4POj7x5L5tGByovU43NoKRbppe
Bbkddb8K1+I3ryT8bnsz/pFaZVSn7QpjSZzZqsUeJDIZsjDCub9zYhptxIIAHoyRLvYo8t+KCMfA
sanbu/t3/0WdRDd4FrIm69XHgbnoqvru6DQHgZue6mmpy+AbRYizvs0nKuo8bJUlfdbMKnGnPVoS
CSYNBDmWO454vm53ogfAGP4dPRPM7rGIyrAwblpp0pPfU4zLjZoDF0QOAkQjwQU8uUVAktlpEi65
soGFCl9SEcaMoytVQPO7+TiYR/lFznN9ZA2A2y24lt+ZmFwUHvy183EAQOyoOc2rGRAQphIXGnUG
v+RVmw6exJKVYsVGww7K6JBmi78NumxfaPlujxTGcQST74yYunkx5EXYo/ArXeahwjeL8M15X6eb
8Th2XOqo2vgvQgofT7OBMDo+BwijShYLPTqUG46PoZtuyYi4A8ZePN12sgeWTuAuMAixMxwxHepz
bICAoL3AIjktuSG9hzvM9W/RhtucX957Ys+EYC1wJzH46hhAspzq+VXwT/+SkohTOxmpwERAUKY2
baJsOMc8abmuzgg2u+ulIAki2iACk1iPTDY3Fpij0jix6d7ePP5nEnIw7kzAROR+nlHoecOp/eK/
v48jJvdM1Pskedw02nXxOEVDFNJ8GxloYrLoqLkJ3LFcsCZvxG/7vHuYXuhgINTkJ2KUrVNkYnht
CixRnXpHFcqjDrL+U3IAtmrGHoKsjAkSnEOxaeQ5WhYCg426XU1irfvQCZSPYXKUHbfe/OkSH0ov
mnGjbGm2yCFEUFsbaN9baRwq9Bbor9T3GPZxw1/UFPAkWuaJ9s5AUXy1j95KrDtOs1x2xjDFcDUk
xSVvLlMVQtKu2eBFd6t2HAOCMPAFkm70dEwohyeJb+iCcTOnaHEA8ACYAn3w9YX60lNC+SBC9gMH
uFfnxDMwhCNCZm+Dau+6ZbgTrE9MHtZhOHP9s2ZBheucyd7+JRS10Xy+lKDTXCybV9wi/1McS3LW
TbjHBR/54yJ9xnxhR4PJr4kQcaYfq3uUkP+W9/T+/yazcob2JYibVTaTMbnQWYEPbW1MXKv4hQyZ
EYk+mEtb2n8cbIvZlnxd838/AAQpFVWcRg06E/0hHua9w8aKpTBb1mErKMk7jy6CD4kcmwCM/HD/
h3xbKi8rblJTk0QhjQs/vqCSmeTs7AUPjOVaByk5akbknEKiVwzMH0A8qFFlwssLUkEkk6/snzwO
q2imI6s9ml9fyMYFkDgjaRMEW7RlxZQnWtXGRsKmI/XOoxxp/gqw9wyQLfz6c2kaE/OgK2S9Fgv1
91g+clvN1BoZRYjBR9v1cjM6SGlrAi43fQed2fZydt9nx/W/zZw1X3HMGuu/Esj6kSQUtGANkag4
MqiX7oCugDEuDBsP68/O4JX8LgdgaZ8zdI9HdGcfdskBac+TZsKUYCVcBDR1c2JHWbdYTkxLoWV8
qntbSrF37jO55VlxmLqqkfaOyi1G54DAVdMV4WSu8lgzkNHF6V9Mc/0S6qhIfxtS74tkC/3Wb+1Z
2sbUHLSpJR3kwEgY5l5gKFFf8AGuH3getRJamJsU7gfyz8004Co43HKVMUnx5UX/Ps4BhsY/s+rW
uOMImDbYpiKWYij9qhCWunHjDr2zS2hW+Y36GM9D7FappFepeqiSZYpKJAR+pXfvQIejCYFgqdo1
24mTjE7QRecBb06wGfQSrLrvB/VrDOknz2ayzFlfGqgLWWeT1LtEYOqoV9JuB23+aC5/Aiezn37m
OBGRhjOSWEvFjrPoVa+OL3VoY/yrGqRY4bDX47ZiMNJSsw28mEcUO6F/bBcp8PRFuJR2Aq0V2EPj
uFe7aogGoQcl+fzmPb6fsUsJY7YXVLz/tj9fVgQjr0brX5PeZhKq7WG1YvOrn5cwZ+MVDcf0jg/E
NDJaisXZSTOxEtCRJ+kykV4BAOGNdMt9cGYHMeUyYmDEtFLsZ6D+7hmF4qhkFgcA3hhzGGbkrMxE
kEVwFNWNuGtjrTQGR//frco7MrS6RNdcvFrC7jrIVXOa/WayWwmwlADnUczIuD3WwyQaBHAWT55R
OATTdaoS3R9uqKRCCVzLt3y3qfKOqp9lEy1LYBPu9eXjsbmIm/Q/sIoKqF5u/iAYmaUosACbaPVi
CmWBf+MqelgRjphZZqZmVMM1txbaPC4kzm2VnE2gMLgWGxWrMg/Wt2NhBekI/qnuV+/UD49OExr+
dEU3LJThmvvvi1dfqG9qjddYSHXeG0aBNp04kgCwcIs+KBB/Mdia8wDbYoxrOwOjBZzZc44aB7Ep
QdVpA9/rxb+5SYhYkGCv4nDynLo1JOh07VoNX0reC+r7S1EBmDamCRqDeGjbSYEvXUPdcuQpNCC+
5qNk2DXLRIg8oDeoISJ75ZVnEMluRv1rqcS36ItLp0pRPy0kH8w/lcQ9dwfEq2YPfo/DUb1DZRl2
qO8diIrLMG4hcrwhvwx4EVuRC4BEedr03pOezv7jLOZcRlEM5dLr4i+2WHjnIurbfZ5wNdWpaNFB
I3wvebiBlRNgBiOrsjRddW/23HpM4ZVDBVRV7+NKI642TnYiqBd2mIKyQjVZ4gd9osbaRArH6uSq
CtDg9jz58LKxwEud3d5elQnvWw6EF9GCLyI9d8CDc/ZqW8QGxGpWHtrMUuVRtmUnn9pLBXe0ZLKe
nDpd6DKyNdADV5J3FxTdGlnFJDKuNaT8h3bLRHw3BPpIUJBko0uAUepwFJuvsTKCk9bOy74pv+bw
16zg4zKQJwLEVjZbK8diMVdlTxvpmTwgpZjN+AgvIBVer73U6CY9QkDtWUYPoa/MgPLL1PEklgUp
fgU98OpUvRY6j2KfhzS3I27iiqscs8zhzLogaUfWTYtEUr9WZhHeoQleU/6YM8e9+dOTkxVU+Df6
HBYX/+Ruj5JmyXzhgbCg07koyRkFhWu6UCsLA/2foffe+Ws4RyLKkXwyqFv2mTV38ah1r0xhhMtN
rXWE2BYqkXimY5tQLGDLVNMf1zkr13NOg1pIflkHkkiyIRA6qBJLvZr/7thMl0BDy4bgUSAL4M6e
YhqS8vGWgktBttBqgyQCH6wXQPQsRnSUby6Aqdo8/ZemIJZabx/Ou39t91zQYejJYKt0Hh0Rgv1m
UdMgroZLrjf4pIIYxT69wPGIaHqezvoCXQgAn0GjgoETPKT1vT7E70Ezfr2+5pcFVivbXbfN7Wwb
pivMfahQe3gIy77AQe3WV8KzIaP4RuYhYfslK/m4hvZtcu/hrmLybb8CiM5PoiGGyl+G0RK2odUs
5i2gkD4W3r+HgAbyxQcCkQRvFDUSW+ymEbxm9cKVARsGxyt5L+OgkwyS5if55BRKmjVrSyUM2hUl
bPfOaWqHGsNqW8tm2PqEv79WmPhkJSoFuNw3a8qBI40+uE+1VX89Gs4xJ5c2JUzBO5JDbj9e7doQ
cSkSkesVmsfkBwoU3xdFu3FyRjuA1K46gSjdY2/Qb2JIeBkVq7UyOv0dCE5Yud+teDXwhMQOBEY4
Rx7vzeei1P2IGb2ZFcE+dkiG2/+FL9pomvhlC/4lFH4iJN/QRSEPsjfoZJT+pPq9zlBH0ZsWJn55
PlIBZ0Ex1YRlIlPUemPXLawlL02UDJ224EwS2Gg+2BfXHJ62veetjtNbmMfctJpVGH3S6gG+Rxm9
Kme5RyVTkFjvBnoVs1BuKQPJVUet3iON1KD0CObBwbH2ddgroXJpOJ9V+55RYbXASSP82aDED8xm
Mdb7jlspt3R15G18Ehx3ymzwdhUcYtT1W2pCTRhr2IK/uZUGVoNTDNY5rFMhrdhWvKRgdmdrYYXH
QGX4PuCVpV9WRY6K73EuLvf+KR15fuPJVyUqH+R25HiionE7mWNajeqtKJysDLweqEKK2hIP5ZKP
kyEitI9baXy/oFR0qIKeQv+PujXWpCw6EYKoLcUPtQk3fy0RggfyJVk+Y5Cqq2cuHWotPtN0gtjh
8cSEKlqx8cH2IQqMFy+hSUHaVhpiT2CJhIbMBlwnwK7Br1ju9FDWAZZu00Iy3442ZW7wO5wnG905
hv+ZP8h9W+CdqxRUyELdcACG3B39ykxrYgNkm2/Diqi6s7EWssMSHbMfEncxQ8hJLEBJo+V2O8Rs
fqiIWklDeBpXDEcdEoYFin9+bF/WdD5EAcwAs2xiex7UwlG0ojL18uKA+jANK1GydQmr6HdoMth6
k29CrmUNdA2yPFpA2Y5Nh5UnFRKuRjxC6XtkHxMYcBEQDgjz4bSpCOXmqfdhgkfAZqSzxxMjX5md
tHprdOMAAqibXFa01sa96emx0X2k/WbkQaIyv/YNKcK5tsvAgN/KlBX/UnlHjRYsNSVWM3sI3J8X
Hv0zRCwN0jiEbRH7QB41iul4ONZu5GLDA/sH4LAPEK04i0f40F87PNrJcnDphLigfrkm2dA8y+Ve
o2xnq1UHVKwn384d9RA+a86cdO4wj9DKU9QiDkQPFnfLZ+Bp6+RiawEdmy/2vBO6nBzgs5rFaox+
cGjzuQ2yxv+oCCG7atbaJ1jMiGjuWuUPGQlW9UBzw/O9Fvhq6089JZnSkLluaAzUZyT2z9mCdOLg
HsQ9ntlpuBORS98IXu39+dSHEWJdEe3G36riit41j5Y6DgX2Apg6JLzoY5HIK6BLqrm95U6RXBCU
6YFjvKLpnDygIEq5Wfc5ZIZPf+xXPub6qnYnvnlSOdVCOewIHDJwBsizNRWEKxgLmJLoyr/raPuG
NzavBtGJpni/YbE/Ta3S8ocxFzspdvJFjkFgzbhc+uYE6du60AIhZpq7B+0xwIzwvGz6pG8xqI7a
mjrqOr/sKx7OEMrxzIfj/4JMtk8L6PTENbzWqUDVceUnn6hnWvWFM8pvOF94FITi/Zy0+AcUhUJf
obyVVXy7f16m6yXFdehUXbf6e/MKs0UwbZA9aQjoebUkbA2fB/qmjfP6TkrjBJ9wqkmZUwMzLfEK
+hTm1Oom/30MPlWI/PyvfLUxzpmWSK4IfN5ZRnLnVwzBBfxxUBhb73ohRwQ36OzLP+p03ghKyZhS
TPysqqmP61GCl/LcSMMF4cgvrZkUTeXhRPAS91eoqI79KS1wnHlTNcFdnVqNZzyvozpIl/XwotXZ
K8m/3YzOPzpw3eLoDa9DW9eJkPI1cPKDIajYwlP2ol8uLllW7QxbPlgi2WpUBMduQRATohLAZjw2
O6xe6X1xPn/ZFrH6e+EhYOtcYIlanQ9tJ8ESFdd8WCeYs9QrT9iKQ8FCTM7UVUqIIeAUYXuFmnZV
zwbSNftw4mrvlHZnwmV/iXmrvgtxJI3eZw8OD3L66TDJT24+JjeezhiMZo6Q28e7iHZLekQk2Ck3
rKYpYJXb0oM50SfRiQ2ZrcX9ZXzbmQ5yy6H/YR66wqR/pm4aSp6VkbWueAlUhYoD5DkZV5tKPbb+
3Wn4aBWyJ+XP/9J8icUzGTDgW4OmE3jZGR8pSsyLTvbJCvquOfgfOQT3mc2ee6m49VaYLNmnS3t+
0j9NQlhWZB4UTevgm0m+83zI2i5VqeBdPcCuO6Nnp9Jl8c5JCLnfspnoplvTRamx4ZbTHY3oIAdQ
qk4vBgBNGrhuScXbVE8+LTxZte/CcELnlQ3h7AVkMJhVgP7W0t/2KPk40CLVdmVgBpWG+YlH1z6i
CxwOTwcmxbj0Y2r9zdfrltN6zLaE4GiEJm7jqnV+6KBi/SpOTZVzQjdR1/6iBGUltyPXcDkRAi6Q
7HfkjoW1WwZoYF5uhnAuuXhcBXSY9avIUNxvPZdS0fxtRUklzxyknYFoP4Ok5+K880pW+KrKDpQu
8r+XDfdu9TXZOE3y5LIPC3qh3l23DqEyzYZe22ZYguQ3hjkwiFnxyL1tdQqKPYBd0zKDNxlKvaeO
12Q2v6VeqNehizlcFsBjLoS5f4V4cYU68DRZzxTE4pEuPjqVp0y1UG7z9gagjEIAIUHQqKAAwviK
yLifWs/+DQJ3TJN+8Ywz2aJNLxgZ/iGnkQ5/9gTdjKoh8A/vBmVAELcoULfilWHKIRv/RNXsDSmV
HHzIWpnhZqXJT+sEa6fJVMuooQQTwqy46fc0ig7uzad1foUh15MCLAGHV2cFrHSRXT54xL//pLQB
BFkOSNghjdEvk9smuYqSxzHyqAVOZ54HoaPoiqwvCXR+C0fCr/KukvnryxCY4EBKCIyDdOt12Juw
CjG0dzhXnmijsVkFNYDjfDf4NqVu3rAQgwLxSz88DIIK85gZhote24yuuqDEWTSWSyqiFr6n8/sH
xSDJfwisntJ/Db6AyeaMFK6oQ5AC1BEtg0Pl8Q7cFlWFzqnHy4z4jm7O9EH7x6XH5e9HPvkSt2xl
Y3CwgS0rzhKyr9Ad2H7kiHGwBJ/7zde4tbRbETGn1akcvPExCYXhOKRqip8Mgb5m1sZOuf7dd+/8
cRgunV9YIIePTEmtN4VSOmMDjw55ADht2s2mh+Y20bekN8D+vMLGiujicC+EgBMEBf4W7s2CZN2+
2NnxqPo6uhronLc1Ow6tPI9uZChX8HVobJEYYMtW6xA4fEbWfBCNxYZcoQ3lMvUuh9vJbr4aZb6b
Eprrd6nDRRDw3yXik9PBWiQiHZ77hYMCmukrI+keiMPHpIyAKK8QQ6dIuWBVtn27YUuxDkpStZCN
ECUQlCtu6kopCvVAyL5zxaquU81Opj3VKeuRUL9MqWZfG9Qt8TshWz7hvjNygOG/3TA6q1LgNWAI
e0T0gNop5OdTAAELpdQTVazBpB4BdRNrHae9YSruR61E4dBcYgfZIW21/v/Mj+dbtmp16IrH4M4E
t3nFJDzfrO53DjQCnE/vYlKje/XgiiAF7wn72MCt/Fxhmxg9jsXTtLW7wPbPhsBBe3O76kKwv3xc
pcq1gsQtatjKrQOd6f50vqVENzuaEyUFNVdIfdcyXSJY07g0ZydvW4NY
`pragma protect end_protected
