`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MXmhAg6x4KfJ5piHHFgE8uACDaO/T4d5WNuRL/TRGDdXNZ17r7ZBwbw4SiFGkk6c
hZR6WQejR0YJUhBq2Lhij4eN1e2bjJilNlkeWn7VolOXgjgsuIlKSh8mkP9mn/L9
CF2ider59YzVQdrZAJIuBR+E7I9n+sSYsRnGu4GX7eQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8912)
unyBfFsy+KbdURyM8innxlIVb9Y6TBHbo0PH9e2zRUmyezkgBp3faF8erT1JtTjo
t+v4ZsZVY4qqZksm2DhDd31N8ZaRWb2YAhNQuWboLzNqaYeI6BNb1OA8o/jwLBn3
PnzCFQ3Kz5MeZraupT2IJKwnXsPQqUmZxnETvV/xjeKhXBu0pLi6Wepc2p4bFaQ4
Zkp6wgYNOwDwq9EbaJmWq5zEGvLAK1YKMbm71fJeb/VXJD+vWx+Y0k1ZrU1ZV6zI
h5UPyOviHiM7tcaecF+rvDUdM3IcN+TA+XZ8v5aSruQAidWVQCh/jxh5f2aUOU+N
yKgwQsOP79mabwe8GSzvgcGjo5m1dVKPEUmeU8NluCDXB3//RBH4rrQja1TxCBIc
W0lOXfOqzmk/DNBMlObyJ56d+o4FrUSTuKGrjJlDcloDXTo7UyRLrf7AQl7ayaQt
IHlKg29AbPs5NrwbCBh61XgfOR1oeJODQbFWiMOcsqrJcFjRETtENBuVc6dQk6h3
B09NcEHhGxKQ334JoT8gGgeM1r3Wkbu8lp4/nUrp/+DlHWR9ZyPNZDhoz8tWvgOh
wQearM9UVsGU1A77ipFjdqy1QsMQwytamMujm/DdshPi+dB6ZpamuIOv+bM0vGBc
Qk/yZ5u+tvlBlVXanMfpW2r80e+8d1qkkUkCDcjyNIQ3ioKf8Gc8NFTD4wuy6mSd
cEMg+PYs9TAHnguTiTy2kcb72mByih/cSBJ18viiH4+qL9u7fayhHrD38qAbJJGz
9ZfMSk05RWeonfD35qvHRgFCaUpBcB66KK6x3qFXzETcB7uaGQTw73dJZPjgWJde
pmwwCxzwudT6hH4ZPaInngejx9UrdBo0wc1H5iJ21m8gVPxcyqBkmcEpUf9Pk/Ns
ab+zb7hGXc3lYslzlxxi6tHk819FuviSMQsa3GZsdCfFP9pM/LBQjFIYaaCtAIUs
DHdYyMr534Jfk5FduOc+bGxDGsY0LJpLV+h6kV0Vq9QV7zUOsXCVKUe6A3AEkfAO
U/P8DN3k6f34HZEYAsteO/YV7yAaU01WwMcuR3q+RmO3gVz0YAdpJJcElHfM1azo
+CXfAeaI6s8ddmlUtPcYXaQQDlKEpYNxYXPBiS7UlQyNrN5rhqdvjjUlB7MBWkiD
At79M0cTkU4VlpUn4jm0X3iUPpFPE3EGzWSL/ih97DG55DM0W11zwUzNW9mif9ub
U2IDhcQkeuSxDHZN2VMIuyaYrVasQbew8SeVOw9CitoJBn3YfNmo5scAnoMFc/qU
SDi0Q8Zgiu6PagfBa+367HraOaG0lXh/MKC60co43qOdoiF7qtOVkXKFbGXkFpTt
BSaBwKFKx/WmZccGChXNiAhyNlmLE1wK0d45USTdhGswHxkJaVnJXVqK+wEWH7wQ
MEUCv9VPSv1bYNQwXwTupdoEFlGvzOiPwIO7YcDGFddOxzc/vfY9vtJ5KEmhFw7R
ptRYohsQ+a8Y4Zl8bkkadVfNX7ETp69M0NtjNw8hz9veLMOkVCir+sQ66hNW6PQG
beQ5UqGizMdNPOQo2Ql3H9UTCgp2xlaHbKlGBFi1kFv6MRvtvWh1BPFpKpWNqQXD
JqGwu5fmIiyGD4ahIypp2bojvlXV1rLr2wBRg5ND0lNlFT+0bPHnxWlt/5KUQpXb
yavOT7Iyu5N1qJdKy+BuIdGkla+wrniLZC/sh1MmvpfLF9xVhes99XhHGfYHxzO5
tPyHXN8LnsqbVT90cJgrhAo1qKZfQyI7oOjk8EvwAUMrE6KWOGybw+zlq5eQdMl9
p/kFPweUM+4vUT/9TRIBSU64CfhHTs9tzcXo6o/tRWJn3SltV3x/P/VQKxH1ufe+
XtXtO57Qf4PNYAU30+6XVRUAscjzc37yQGDagFay5rfmGTkEFnfp+hpjzs058W8j
QUsfBBhXUmWvojyFHB93OIiYP/qtNhS9/S5hGpobbFW22h/an8WJhq/1/tWeFU6D
/t1rPqlJoChwjnKiXRi9wsLMabE6VDLGPDhHSzdAp66cORtk0sKuj0HfKRkill67
yQ89jwNcImM1LsrzlFlVbDcBsoQBgi2d2Xk6TJzJNfzIrF5P6Lo8B42n3AURHypu
JD3UPMUcb+f2wZxyEYKH8TRPwgCzp53CoqQg8vasX++Y2cmi7EUR/qxiGdT6/A3G
V3rM+CThJ3by5gvbH/q8ENqZPzwcM4qJEd7uJpLsLcBzS52+vE+dBnDWC6T/q0+Y
FtStJ4TT8Tc2Lt9QnEU/hQ/3he4/RioECtjjVbgvVzOvI9KRwHzRGspZQXiNj9D1
4hhFMpEghwfYV5dt2+TTKdIiGd93WDIxAp6oRrbi1UVc89IJ4SWsxRDPcJRRMxQJ
9nT/R90j8vmpkUH2FSwR6mQnxhQi/H8KtxHC0pSnLwsESYaL52hG45+mKsGjZK9w
Jh37P0z1k5ZtFYWmz6VoAMtJVdkXyy5NFoq/U3GtDzr3iU+0cmM+vxQM+NJwtmo0
vxLTBKPAvUj3w0Muf8LfqP6KrNMp9WR8cB/9mACoZE2DlNy/nP6OpSGWEoNm32jj
cWVmKQ3soE/DrKbdgPG9mjbgz+4G75Te2lPatoVflp97e3JE8ghaUqqO0PKAEHhG
BEtSZpd4cSUizWaUqa+ab38B+nKoKoL2ntuKqOuDGtmk1jeb7F76wCE7xFtjVI+R
LxuCnVyqCKVvcvHlwMJ7bdXlWnajf+87k3m53sXvW6vM3NDd1gcTRAjaPKiuB14R
SW5OPicojV4wWvyRjwwGaxjOsikfedGjsZEFSoQ7M8ojJ2nP43nCcgYQr8Msd+o9
0UrqIYSeBNw07xxr7dbeg5H/gvraaqykl23sTKPgsqYLOlCzvh7zzXRHNIpYAobZ
fw4pVxQQLnTL+7dJDVaob1aNXqTnCC3XCsrW47X1DscPAuOsJnWtB27uXWuaJlgy
8SmK8/TfRcq1OcRF6Foqx/vTRh9CJWGBcKUVLM15mv6aTG8OAVqq09YK6Ck3kCul
B2EEPKm93DQ5f4gLOvXW+02yUyUlIEZ3jFCPsS/rlzHHTt7CzH4as/OqHaPVzFkw
XP858dxbBxBkRDqMMClJmubp3hGtNYV4odQz7z75oT/JhivEDCHCNCvNH+3yx5jK
B/tHxNUXYmdiHcypEMTq2GEHRIHvNioa6ebgCFRuAwJ5wGnhVcTWeCiPvKtLLLe5
6UzGzq4J/W358r9pkYgw4t2+HrckiIUkU3NZgs+1RYYKWMTSzljrzzyApHoW4TCl
c8URrBQX4rWC1JkSaPIczHNTQNxiUyzgHsOfC/VzhURqZw00Uie+SRnQaZwNaZzO
qIbPftjTQcSjimE+bMq4suJeGoUFkshATcACPgW7zwsC9bXroWslrz11eFkQQhAx
u00I9i8tiqMSru5kHB5J+4kEPuGIsWfF/0Q/VHJMLfQUziSDM/i7FrZmH4y7UV44
hSPdgF8VVCxmRa7+TNhEWqULuCpDobZDM2g85B8dTpiuBH+1WQ5F+FC5mc0uEww4
Rl/UAcRBgiRWKraKrSudSdj7okG8tpWLq/LXem1xGc79OL/HN03dUJ5+TqVowE0q
zfE6VGXfHr+Sct9MC3YLmccev06kKhz8hkaVAadRab4eV+n4peIu5VUXIBbBkdL6
dj9E1MQtxNqFrgDOjZI1io1xyuNvbmgOyEmM+7O6FCUdqf3siFR+MOv6m39VvWJ4
92y6OonQ3qZJyrm5pSokpcGz0zbrMKjoORp5AEdXYiHu+Xbkf/rQTwVAx/4ZmaPv
ed89kE4+hSwjB8Rc/HTh4vj9q0Rca+b3QT0IrwIE7RTkrod8j9C88NL66QsPbxhC
yn5reYfYo/FMBeoYuuaKTOK5s7SK0/ce10OhGtLtoIOZICLMNjTypH4Nd91wDQ5z
C4GRBEaXVDE/oASN1aEmYYlftLGLIbcwsvMMDOFU6uEQVXNPWMIvHA25Wm9z++Ia
OFB9EaD8sCKO0NUMm9XvKdpFxNEAFrLA0KkMORy2jEdRKWoDicBVjKmYQNlMj/7Z
cEOG1nedBOJydT1StFfIs7xVXeK8PU48X/cp2xUEMMzc0IXOSfknsKk7bxa8ZouF
EcsUDcJJC+ib+kOabzDaNCvguW9rc6I9k//mO5643YwjGl+Gh+xzXTO9NIv11oSw
1bVHWr1y/mlvGOx+xNVmVKYhpOOjZuaorEZpyTCopgDjw4v5DGte6Gz8i2ggw54N
7P6gKVX1uWSy8kJMeVb+wGvc8R3ZRVJg8WKYbXl91oVsBu/abl76JE8Ho0wAn5Lw
aeQNuqlrR3WdVXSTWXgkghqge4ylXnKIq29k9mANJe7n8h5JA8yArkXU2a8C700u
H5TZqfj/JCJsF6OLpNEo+QiXlhAS4nckGD84DXTIFJlmOLHBMhfsREbCgIv9VGM8
UaJSX2uZS6rN+o3XUDcxMXrQhPbTV4MvO6PyuDlsKaYjcyV25QKBy7kWNkVwrhDz
88nCP3oEbLZYEorVgECxMXDBbSNt+lsfJN2A4Nm0CN+ypzUWl/EoKgLzFcDe/QzK
0MYLE7zfIJdns2W5i1EP+lAbyDgo4Qi/ApP6UW01rGgE8o3pi7tZS+mL9X7PSOdZ
MD+alhmoje+oFa8/NdxuR47+PCD1ghFvOCp3qc4kAhGSmz6Qcj68mduD2ExEMeki
iIVVKhBj1RF63bCkOHs4k8Kk/xBW5kmh/lUxj0KS+r2o7OrxQubsEvuFpVcPWAVl
3wVk5c0N6o1Qx1AaZQRQmN35MkZeRJvFpXg8gVAPbnI7KyT2SNU/FBTijrPiwDTr
d21OjbZd+l7CjMTvIBFMxF+Q5mTGXuGxinwN0DeuhUWq0nhsi+dOT3G3aLFrSVyM
88WS+Nzd1HV7pJ1HcnMc8YvqoPfJbyc83mMH0AWZJt8wdsscp8GE3wi8lrhmtTjb
VbpUyKwvhdFHKs/dfvHjA1Oh+iRiQX4UvQrcIfKvG48WGDevBJD/BEFJRQuqbvUM
ch549T1C695xhgYh/VVcfboUlaKENhTMB0nRPenklfz+u5DdGWWnbKOOZgah3wgG
VU2hZQeXZBx+tp6t0NZhh9icodO9A3ShhUMFb4igc1+a/XvZIMZDvNPH0J2PWfEW
zGn0VgKS4zBXr++pmLraOTmlGJsLkhYO7xwEu+3dluN0+h4mO+NyfAPuKlLAfM58
P2dR4EHaB4WnseL+UKMmQJofamPAhbc4fJZnVoJ2X5tbtmNHT/Kmp2qHfro8gPK5
ZPoMMDACmw+j3pjwrjh1Qa4NiLpm17SEwwH4xQiEdUQDnmewJAAHB0tHjUL/1sIM
LfJcV5YI2+gR4P3E+oGN9bFs/dTIs5nZxwsyNpoNBdq1RAZyAgkXDAihFwAnCRNn
IKyjineQAMs/tJd1/hvWvrAmMWZmdq4EBqhXRvRYz/Z2plX7WdFsyJO5LxV8oBg8
JG8GXr4J+EyIPmifMmGoBixOZO3Pu74gU1B3EdiLfRqJAGdyrjoJyfAj969MobS2
B5X06RCaAJ7Ja7QK1ASx0uXMx6OHTLUPuVk96pw1fAOI4DPP5Edwdxc+iSupFctm
XLrgE2Cw1jo8nwNcMHFINsz0Y99Rt7uJStf6Qax/8A8g07onNufBgXXhxIeCpT39
K0LiTUCRVPhOCuz9+SO1CxDDXqPgfCcvLkdVHATGmJ8ZxmUlwaCj9er+IqPVC291
Z/X2tXYaSNyqqjigc5baoD9E7cpzTikZ4aKQuRi7wvxsIojGKJ4rIebmNLJYUjSH
qrHaewzwAL8PsjgvYpX663LL9fF+7BZODeoMYG7FTKHjf4pTfiZaKG5duw/TfORy
+OCiCT4x0JU9ct3wHGuFnhyRJNZUblRDeqxP8Wr2xdFoJgWOowOxVZn0mrWsSUcB
HZ6z4g3MU5z/YCdqzFXfoVvjGoXuvjk/3CQhwGWO3h+z4UB7D9O/4zse/kF2Y2ce
4N4cc+G83zB0vdUH0E76/1LMhP/ieZGIvJ8jEcns1LsUfZcoRSDKU+UZtPbzOL+5
UAwfowOmIuoDpjIC19lhjKu5VAZF5F6nz6U7TC4K0zabkhXOyt3we1pxedfyF0NC
qbLp9S+b1ksTNEe3lthJs5yPXF1zOvymM/nk13PRtMvzrLCHVfA6gLRRz5SLt4a5
okhekk8+pKW8PfO0bGdYdTpMfWX2HE6SbaM9mSbypoJyMsluXkidmYWRN9BaBzDQ
Jaae8LjWsTkTK74MmqebhvwSOcITTNFyPLAWt8jVzGad7RiT7cshhdLYRkDGxkFe
1VPcp7riM/CZw0JhGg4+iaeh+PoQ68PcjLTDXLGn+xqFIO/4yBh5dHXkLGxPTpiX
VZdvMGrrcFw92kKwPbz/eLHiUmH3mpCrKwqqQvH1671FFPd1hUFZewBVnm5xVlbE
uaM2t0QAldT1yTKZK5lJUGJRyV7XI9Q8ATEPS17N9JE8jig/SLUNvkLstFy+RvCg
gUKS+CBzKdHXb6BK297dq38i9452sjwo47At8JWgSkuubL/CHkJbEKSk6CVZpm1T
w2ZEhksihERIaxEK+nJ3jMvlTPCJWaY+6pxNhyauo1klsaS0tRSPUHLU6KTc4jbG
btLnBQQrjslCcCFovVUmiE+gjOTJq5D2zzdNMyel67WGmA6VemuPgQ0dfFe5n3Q8
9rrq6AVhY2tH7w/XQoQVW9g75ZZ2XIu29tS7PQPgDzya77BdsVf6cAuHYHUx6SHE
IWorXqLw+cGp7oRgYENpIZ+NLFFBZ0oS+lEfl4FxxaDakETQCdbogBnhBlLnA2iK
3QKE8Kn21GR3GyU6ZE0tJ1Q0jgkNcXvqry1jEwvvQJsExFdOfhLwt8XbRBaF5rIW
Y1ARxmQZt0iyMQxB+eHoTur1PJAfhOytneF8+EbOOCEP/+PpkHHYos8/F9Y6OJpL
S553Lju513jdE9/K24fN9yMTiXdZXsFDXWvYMIQeuGVdzDpX8tpRNbDv4qxH+EBX
qa6nevFHVQUVpFtfNP+pJ0mmn05zEEAtmJvdGdD7Y63nlI+A497fLm/OvHSWI8NN
UERgiM2/FjnXB4UhvWkgxLlL/nVX8InzbzbYVvGd8zt6MCo/Z0iqz8CNU6bSbGI7
wWaCk5/LqjN3WTHiCxRRMBY6PtH1eo8mFGL0wlnsETgHemUSATax6RGvl9KvzqWC
wzHSZBgfN62v709UVkLUGwnTNxFynvAbyxbMneKygtTRLfx30YnnmlDsIrfPlUxF
RPsHTlNvbotspL1U5Tk4JufAQGysqqEyydu8zvXfNEZYcX2TtFSPBi7La3g0/ith
XADDqHNiBa+tIYSer00uxHlyxVUiVkXUp0qLCLtK2KH3htDQ5yqlcprez51PwLZl
OlMjrssZd369zUUkVFXYBfSxSorv0Ch9S/YOS6CHQG/3REqXpe6Iibvr77Vl6RfA
nFZJ7YP5H7WQTZa/NKiq6uN0ilAQYj2mt+UL3NsrHRpx/HkToqP0Yz67dvVnnXRn
aSG47aV9ygszZcqougJhlqpmjZeHYuAFFMOh7eRLaH7CGT4pXpZ4smjTADif83zT
njO6ml4eh/J4KcwWuHm0kDoHYFx75pVcZOv2H91zUtqgofHz9YeCjHHgwfBe9OTY
k746Hq8drrR0Tp6Oq1+bemFoUEKw+zsjKd7wXq9BrwB67QLf5blxQDqEoaagJOKi
ceiZ/ArPOzSL43j6kEO94w4aEdrneVqWvwHMJAPgVRVfSG1SnUVPUA4bCF0xIdPp
6KNx1PrJlgmgttPXTzkIumvVKkyTx0SmctQ2AvARSZ4rreYBrfr9jzjndz53AqEG
p03pzdxUcxKhauwaq9tMfVCHndSbOCcacKRY55MOK69/oH6yZmrsFMR7FWKVcByH
s6cDLa2kiq5Tqh2AZcNsPz96u/UL7YHAgiWIhhd9SVGWDUzijWkTZ+U/joX0vqVs
y+uaJQQhoWAYrJvgc+dmCwRD6KNaV0O1FMrMnMuXZASYCAw4DOJEX6Sv6TJup7nU
REuKueZSwCYrzEicjeJjJqOyz2kzAOUgYrJqgMzvORInP7IBq6hZJ23tIGqzHSuJ
OqVb5uQYReokPUfU3lL7JHrf29viwry7Xru/9HFPEOtBZ6fwLOARW7fSJtI1oWqV
0HBdfiGXip6XomqF6lwwayIX3eHzoq64yw7tqmF0ir6RAoeEIMQD/Mv1OYyAnzCg
/QlOr6fXhm3GkwqadfEzwYBMQaxpKcBVIdfHfe2SDqcGFjBM3oDGFpwLUa4zHFdY
vWzNUhiBJ3g6f8p1BjD91Jq0EETlhboIWmRkMGIDrsjz9ItpU+kIGqctr2Ce+kB7
QSPSmwbvnyDb2Ht/iwlx2QOz2Gs/fBtbfaS5wNYwj8YNKqIjEXITLbIAysXpboLx
G0K15k9EpLCTjJfojcUphQZ32I1gkpAmOpQ1dMNRNr0YHsmKge9AHvBsTHMvQKQo
OePTgZhjNlIIL73RM084+6B+W2I3mMbybgpAjsGJiNN0XFrH73fSqTL/xTR+kdOn
p+iXB9tx5SA9fSYpJlu6lWx98d3X1JKfZvQ86fP4aND6j6PAHUK5Ns8Megl6qb0C
maqO4flwWTEoelRbnAExueV95AUhj5TMN86DJMtTKgc6adVj/OqoiJgYRxDCptDv
zIxzOHSTuw4UNvdfxIUCz8qBPZZYbs22M1oCazr199vXmPGmUO0bx6JW8fEoy2ko
SuwLRpevDb5VXz6kZSrFaldIDbd7RQVMEgD2JmCAiBB9YSQ97lNlgmfkIDrsIRMR
Px/qXTc26kRdjP0FFk2VISgIV63mQc9wkQtvNTesRYCXe24k+SyXrFBb3zuOYHKs
/mkAbR2/c2TsMSdSCe92P/hCZjnwhmunH9hs/xHjdW/2XYALHtojyoPKhX0qJicq
D8vWN2O0xiyc1222I30NpDYXOTjnlBarkVMwyAzGZolbFfSDOyFrH0ETF7xcLMWl
ZmHB79flt8x090985ZNo5zVSy+Fndv3c7Hm+HK3HFe6l9rF/wiQFKY57ACnZnOAD
RrIleRx0TnFyFRs99Zov2wcgf4nQWrUMbaPJG6B/8aGAiB6otBPC7Pn4ISOayLRF
iNLO7wGx3pJ7Q9e0S4Be93KaM+DnJvj3Ap2FiugxXSRdUTKQ90lQKE1c5BeFouX6
wl6YnPpabmqYifwoJK41+BLMxG9o5bKOi0STNir0nX2225FF9CPvByBTrZZT34BI
vgGT5u71iDHYHkVCYP351IK3zW2IQcVMt5KYXKmDQM2/6EsQS7gfozcG6rpym3t2
g143WyEmTDyHi4zxZhF9+VIRv9l4niHrirzFnAv7NY02BhVnuKKhPPbu0BBXUlnM
qf1Fbfal5RbY2SiuznTM2JFGPkPfWVwGpoR6lyL/00GjNN9rc6tpZ70aCEpu5xDD
BEDauwjJehEp/QzGYYZm/cp/KoWMefLfMNWn5/gsKf3Ho9A871poPp1zVcT6rlZN
RD7bJO9+myN1il4Tk7aMG938KDMmc5o/61Ay6xgSD4l4YydWbjjEGzN7jT9L8zKQ
GC1SPah0IpXmBr0l8sr2ovo1N177ECLqqwFdRY+hukfrxw2t1/5WZC/X9Bjt07Li
dOFDIrrjRN/trTWTGZrczFFi0hK8bQoUIoB48Li+lmRAm1wU5QJ7EuA178ggnSw0
I43RM7RhBG0d+Z5EoqV0ttjRyWqIfPd2qPggyGLOgq6GX51/72RZemLpsg/JqCMO
YicI7cSTA/EOx2S0TEFB9QEWgFqI9yKv4rd5CitHMSVexvPmOcmV0IcuhnLtrl6z
aZxXD4CyhIv5M11BXjsG2/DapgXr/ucP8EbUO1pTuQGDTAomVGT85rYjVAING9ft
tps9DkviF3je4PLc1Xj7EXGvEoQjweHzPJNrVuVmNqarOuU5oEZdm/d4k2YLReqi
sf7BNNcpcORnRzw+DkPWHVO/NeETVb5yVWEgEA/4Nf8NM5RZ6B7Vq4c4jhmgQE3U
YY0qn5OsA9Fqogcrw0vp7stDG5DExkiSkHpq2hhI8XU1d/on67ZJ6t62se9ZkJje
rylLVaHvFmx/0IE+PoTG4ga0W88JqWAOO7+xtv0JeSpWW1V7e6sq8fzFFSE3eBZP
LGJIvkvIvDZceC7iRakQJ3pL8iRCPVD6m8wmk19jkBZl10n5aO/85ckOkDc0BHL7
WSd7kiiv6d83rr73f8AAQD+ejNmWRX4Dxqp26Jkepr/Wa9Qgb8y2xEcSWSL4fmoQ
35KcH+83KgtQba5W2GM9ZYY0C2vi9/Fw1ApqZlzv3l+WKFh1KE+YYpGH+VGFugWm
hoxCPAu07BhLNnd1zOEgzw5OTe20NhALfP5srBIMxYJeMIupXpUfChu4FQqMXpmT
7y0XhtA7+c+IteGjqsPkV9f8fmF23FzTrBEmrj/yqyYaiZqdSsEmgSUA0tUO7Ibx
IqMbvruODn7yU87VbrY+F21a/61D2AJSBMWdiltgqli3oabM7u8p0MD/wDOujor8
7I7JDBwdibQ6hWCdpEKtxqI5vlenqB3GfKKbqey0JEfdvBlgBy2Sq5+0+deR+GRi
YiOppwBzih7O5Dyj6O1vpXqOr2VEh9J5aU5MaLK0xuxM+WpE/wKjmGXIEm1ppM+8
QFSVBw8olAGzzMO9YhTuiwKgWJxtwPuBguAFpxuifl/yj11Pc4ADNPnApXKOtucH
AnG6dPTTTCuxCKfDl7Vmx5rwcdg8pzQnM9IhWg41o4IfnLE2UiN8LfO5tu8/06ho
0bo4Y2woLUlZJNQS4q+CZERTqY4ZvOOO2GMR6W1j0RRy+37lSRMyuzVKmds8XiA/
tnnz4uaTPVL6w6NxGep+J9Sfo/9OwlF4vnQIPhCCU2kYaMPQWmlmy9xlvAU4IWfg
Ko8WSwbKQXZX5q1IN8+y3d05+j2vJMMABNsZq9PDGi1RqvxKgoo8bsP1giirM9HQ
l+1CkZ523UahmFBH4BwF7YHCyCiOOehpIDMZ0Y7odwqC6oKQBJuj7RXw/uAlFTYc
XupX2WvkvWn5aUTJoVEpa124aPe6I5W0xCO9ByUurrMlK17jDbLKA8P8pIR0IboF
69mhUxC6MfiIHCIdpLKRKqIOeEb75h/KXmUyrleAGiAMROLPq0ROYJHWTvbi3CZD
AIw+S3L2wXZxoc349OfG3NwislJZHA5zoHjUTS+cocTUvsv+aPbfWM3EEb2JuzXr
i7truf2yq3Rfe7ra/ojcdfc8zJBqIGn96AUT7B6oSDr26GZ0tI78BwC88fIgv0de
Na1JWohsHYnF+vlrPRNBwgNF0qXcKia5LN+ipiNNbKkbLAoAyEeNb8quJAjt/Pai
4QIbLGKkRDZCEPKAK7OVVO/FZjffwKAxqRZxZJ9fob9TWRYyeinh3WTyuLawTD4/
OMssxMuCUTGUI6phDIjlld50cyWYYP9sEwDwYFQXTpIg4rpm7qeAj2/MKeyXTJNF
8QaQYhSnADDXKANVwgij7NMOBJeJG84WVji86kec2nXS1oplnBifIK02weFyB4ry
+mhSYuPJopHqBJpeVF1u7YiW6wIMDlGtF8lZtuINBZBnniXDeJS+XvtumpVDnjqH
O6PTMKX2syPRbZo0BviHnE+hEY0cIjc1wACc2SLjVB0h6fXQWrQPINa0j3o9VXik
RQgl6cZeIn7wGMxesAERx37xqkNeYFF9CBDjJ7FYqrxx7nn+wpxezy+WI2EPMmwI
fPM7ONSi2PFYroY+rzZ2GouhJ/DDqKQ0yJ7+kYdYvJTF4OWNG6x+yfIKSTlGTiMK
RuIHYmhlDzBoSDthf5b7XRka14BlE3807Ohrdqf+bcujxtB9C6c3JOTsvOQPfCBy
ra2Zz6Zyhk5S6ca9O0X4F/1j9HrtCWSC8sLHe0Uegfs=
`pragma protect end_protected
