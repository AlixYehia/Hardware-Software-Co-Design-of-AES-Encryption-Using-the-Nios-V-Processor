// AES_encrypt_tb.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module AES_encrypt_tb (
	);

	wire    aes_encrypt_inst_clk_bfm_clk_clk; // AES_encrypt_inst_clk_bfm:clk -> AES_encrypt_inst:clk_clk

	AES_encrypt aes_encrypt_inst (
		.clk_clk (aes_encrypt_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) aes_encrypt_inst_clk_bfm (
		.clk (aes_encrypt_inst_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
