`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VyhJRrHpTPWCoApj1htLxaAYbbOcSyYQr1buYlWA258xmV43aUjuGvdXaLFvO/eO
ASNJuOIa43UG7ShtYr6WSavGbVTHkbb4xhHlnv9cPH9zFclZBaKewWFUCHpssRdw
KHNMTT4SAMMCxclpd0yv64QNdmxiT2+iddK8l2d8Vu8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9520)
0EdVrb5mQx0T29bX+JGQ3Df0bSgFL4unfe4W3Y7OW0wH8zBHWlBjDp4C5RfGcMsa
CjkAEvcffyLKQ+ykJaZQAq5IFVaZ5t1SKuYEm3dOw6iI9tmrwDKN0gv1gGNy2a6S
LExkPngt/u02eupS8ZKP8oVYK4H11enTK4kkh+r+RHHwInh2oE+1IxDSmTCMm+pF
Qil5B0ax5hNRDlaqaCLGcizMz0T+QPdShpPqxABz+zLBV3wh23mn3+mVLikfqu9s
TIvavtFm632lnS+fKRdgmaD4hkqyhcOTjur/VDXYUWxbKyJnIfQB0jh04IPGUKpy
x1QHiA1tPka1NZlNZpVxi92gABP0UCQrMA9xfilfuQg10MaX0kI2l13FjYp+Fh31
kQ/t12OyVA+gYzFXUgLrQPR2fhOw57GzpTkyWvcYIVKCuXfDbC4j4Plei1gVPQ6c
uBZOiyHbhpIaJsIvWVirsqjP3I1CPvZ/UP7RH1qJspSqlXD7ZwrGXkhk/RyMjTOv
5MOjOKeBkXxgrmJppm525Mizcs7Rd2Eo2m2DZWxAvYcK2Ny02gHgfbThk6Ncbnwx
bfLJXkRWYHCvtYgCp810WmJSnbP7R+Ti58XxlnkgjfB8t34SCRDDwbRx/egKQL7S
oR2iJYNabdd0k9FoWgHYOnqQjGFdJ2WhHWu7PI5axhj3bksuI09VkYVbROju5p8D
hKFgDB7bo/2OZbTfirWZWzuZ5pD+YBaC0kVE962Uiw79FqUCFdcu5siKFUSknYTv
gkeDn4X5dyc5rOIS7Q97EgE6BRifG4GQePZ6roKxf+3+FslmIQlQJkHU9+OGz+1g
2Iw7vTE4vcIuOn3oQCR0ezwmTfPuqhiAXfGTyTsKpMXF8Te6VyT8X7ng8vWX+MiJ
kuWmQE9kxr6FhfGCLYeSc96TvMdZKT769aLt5TcAbO93UT4FcEh4JMsgL4BQY9YB
sbG+jFatp+RZ3KLO3N8xSXXqJ763DF4JOL0fBnBIHcaxPCKsoK5ZVmfM7BnIM48n
8GMVDLWhfPbcnKR0xetk+GAK6lw40RbdVts8T2X6ZA/763mWvy6vr+KSn4kpQoIz
0XPiXpywyFi4nBttSSkCqRawwVO2YNFV7HD3OTh1Crbkif2UE090ejd+HRc2f7A9
WZUaibnaMSwl6HOPMsygmhai6Gm7azvj11nwPsa/orFIOou7y2uw7HyEAuvVP+W7
K/wMKKu1/51m6PUJGDP7sGo24gp81OPKtUMpEjyd82Oto1F7Anwcy9QeNVOvVT+/
GtTXgXGMH3xvVEExOw+iYPQZpjD6OoR2+DmMdBD4QN7IO94i5+SpPJ9U8S+jO6lt
AYfJ8ZYECjEB/O1/bxPd+rUCjlMhG+UTQvLfRlGKb2/bbnVNPAVP8MUigcTixI3p
BLRZ3hjOzl9447gHqU0xf67/j+NqHO17imUnbN9VAoN1GVimUpGbX9BuGelFrFMY
lGuEZR6y++1E0Ajvj6HboIhv74nBzoTn8GNiEnCwRdhQlPc91optfEfBMtuhVARj
HLflLawFRgcVphxjxExFgoU81ur8uQU7YAj+Kb5Fsi+/gkD44T0DqsdHcFQlia6j
Uhkkrf3pp6VTmTOEqKk0nBwVARgYwrWavEB2YV76OgiT0gFp2O2W+zlAW/5Xr7IO
k7YN+ewTa0z05kp18CuZJZ2O2HJzlbIcXVffTkWUq8GQov5rrdxGunFqEumqz9dR
KWas1IrTP7Jo4QbyV9XKGhU0h2Bt0/LoUJgVF7Pm/JAB34fkaO4P+ogHZIL8phTm
gbshW0jPxBeECTcD8rWXFSOaSUrrRuDAVXVEY3hLgwhZz+/5ktVf9Qut4uSeC8s/
WiBlGKsGINB0R2zNb32rYCRoDIuzhSTyDzhWoG78XhAi+sy7SLRMgFIyAVvxbqE5
jlRdSpLbaal/AONv/6iBbNMdY8wUKMnbrLavdBH3S5B5tpBGVNZK21KHFcyMEWko
3biJFiTG7+kz05UDUj5++SF7+BAVH+SXKoHsdJVbRYBXI4SOZ7IJsYnQrc61MoSm
R7wUDh9ROR3x3y3fg+NxuNDEUJ66OmERF7D151VgcRAlHuCiqGNUgttUkH8LO5TZ
wN3ryciwj4/+jeXOSWhfO5CvR9s6v1puHrFDxi8B5EPUjtxWuC9eplKL3AEKRlKa
JSggqHoXDo5SDI515eksJvzdwcQjnTkokpa2HAMQnma50I6a6QFwAHrhf0kXnJu/
ouCC6Ur4LdTjbJXuTDZ+9p/vIuAhzvSDYcmIMQXDX2uknf86BDNA1sh8/FNi+lFV
T5tOjvp2/XACg5Pg79+8dtBlNEcc1opSttv6Igch6ljqMftxtFAAkVvum6KSpcgw
vkMs1TQ6ElRv2sg/MH0WlR+HiYAai5zI1tmPM5tPbc/e5G5l9DWHiMaFE6EDGMGg
QWCfLvkaTNQj4IQZoZfR8YvAg1Obw+dpYUoGiNwmsWnMSsiYIA/R0FS/GASzrDTU
Uqaf3yKByS/nW6SJinf5ETYZtVDo5dZoQg1Eb2FZBgQ5gZpXfKYuDDJgkuxleGfB
+chWhpnxDpRJsnz2+0+b+PtgPE+voo+ai1Wu2L83KeuyXkztAjT6LttndjgaakLL
x4ExthtMz/l+SmGVGbvD6M1Yh7xI1xsVd8Huam75izPN79RZFff68i+JZ3fhHHaR
/t9l2w89w70TTwT72HqG8vExxG4LLOatnY3uAa7gVF2oVPf2yv9FXPYMhxEHcEDb
ogIn4RSKI6XyvYxDSapx3pxBSKMz1/NBNDZtuDLR4ZPRbSUQrh4pW4NHtGEVGwVH
i0HG78F11KMOeZNS8sDXR5snUoWUiIxlgxq1vlJ3Raxa2EO1ElPPz3Td79hiwXcB
qxmmuDFSI5Q81PIsmecZ4nypzubN09KP9dfUR+wkZ9JMTQmIOWIPmiZ9/Ycxp1QA
IO3PZs2Uqr5KlrXMH++90FGENwG5j+ybiLAHDoHDHUT3xCHWoBlG+HBfSp0+Fvwh
F6uaThL4RyVK6sax72ydnJniz2edsbOhlOu2v+VROclEqcIIH1mX4H92mUyCyO34
xHJlzLPyHfEMKxIELE11vxHqtWF/3XCHGOJ3BFKmFFjO/Ai/1btwHmWevPeC/0nC
bO3EPVbAQvM6eTwRIwibqs1GM+2FHb7W1+OZoVS4vJAfwWw1M/sz0IAMWdLj57Mr
RBRrcVDsoi8+fzEmZ1gn3B+AxNq3szk4w0WcQRMEXoyjZpbPboQMA4WqZvgexNqe
grFAO0ZctOt8qOq8oM+uAHj56VdtSThoZk33qzPWFTGRMMO7R7uj1lkcRHdgEmsc
7dSJacw2U8iLtkBPp1aN6wVpkxLSy9+saWMcY3WMngI9EzaO5tmpopdPQcQnCLcd
TK+VtzH9X/UcAo/PTnLBARiW/2Tvd8P4T1mJybcFRMnzFhyPySg6ph1UE3oU5c00
zothyY6l6sAauZjmfA4P4ZmXqgxmZmlGmIY/ceqXPYMu3soEaxxze3dFxw7mmQxP
+RnMf7gl6pxlE+VCPAJy1IBHD70rtCdVbR+LzpFkS1NR9czN7YiYJ0FlLZTSikb8
QpfLdOp3eh4in5gxUt/qyrKv+k+WtIDsUkL2SnHihNrbbw4jHxkxQU8p4VRh3vGl
EVHC3F0ipiPw1VXFey3zJE7sCAl+Kpmph5IWreiTl5yeIgnY4epaBJHUCUj2Ud95
HvqFuBURUQZlvTJP9q5iXcpDfyieZ6aT7z91lNvulNX2JDl1tMnbcTpC1087s8pw
w+aq/RisGdkNbZqzAuvK9AcgPwmPebg8dGWyLTLeZCZQTK7B10DCdBZgBhHUz5nL
u0l7jcWspE02Y6+knqruKrPFCKDLIzz2q1Ub4V1Lc47iBCP9Wp5vWZOCJjT2/s8S
0RFwDJ/geLjbnBWtocD+dovUQlMmjRtvKTs6U9Vee0lAYDLQ87k1jbxbx9xeSij9
uGoMrtsXcQI0xeYhqkLo0w+1NqIBNefzUOnHLzfLPZg2OQFx3TxuW3fzAForaeBP
mTa+XDham+iSYR5QerhmN1YZIMd1vYBahX42vLu/yiKKmNhdi2fhbeDH9ZPAUh+N
CNcWxaWBOkziaKVqGKcoZZXtErhNejKGfhwEuSbw5cQGVSiMC1uea2s9EtsgrZWd
lZ/KYpqlSYAXnBtm9KAXOo+dmXXgdbKm7bH6wqhCIFDH/7rZ+oDc2fU+0fopKN6g
HPrxywYlgWA/4s9YquJi7K/MDCKF0BqZ+jrNNztIZrtmdhOnk8pK0kQAtGH4pjlW
Yy+zXGKQ9v5lxz824UrdRZfqrQO5+GcT5gJ8KI9TzicxQ7jZQO1JUkqTcS0Frsmk
0z/dzOCJvv2s8BwqUvx4m7YgUIrSV3ErHVx9bPFtx5RrKRG9psxGQLDzLzH4xUj9
JGxA+TCfnw5M05fR1mUQ0vfUIHB4+68ev61zwQB+3x9Y2emEXV1F+EJUNmj5J4Md
YsHNqY4IN+kEqMKGIrNUfvtKyJndxTasJ1vceIlvKUxL3krZUqkI1A7SFdbc4atB
zpXkGNYXgmwRWTp/Q5qL2t668fAbY9NTppc99VolSohP6QackeBzfixodYWKbjaw
aD7lmFONomGth5QCQcJo0tbalyUmIHONDU2KSma+RuFqM+GbGX/Yx0UCF7Zyzv85
5EsNHKkqGlVj4fFYETUQlkBM+TKxGPLuqummmst9IMONHO7Bnn9yeZMUI52OrZXY
UYgy3SzuUIVsfuSV1dA46vrzPm0oCnM9ZSuAsfTr3txBGco+TZukcsloTO/zhCqd
RxP0HEEjfdjUbwBS4KZIP1FU8dFOUp1W4qKcfYGfFCbEbqMJbDGS+D81Zt1jqCLu
6J7DrYywgjnRQuCbDSSRR8CEE/1PzXJtR3t3uAjyXcjeV/vzKDTeB+mmZCoHEsvB
FoOAhOVXnbQX8uVN+yHBzUTQe1CXWvl52s8vIE/rgg7GVO3sR9G4Mc9/cgiXifoq
thwQ5ZSy9c+cIhyFHoMcip0Cw8KQOfNvtw49izfg4BPbkfcVL11O+QVBtewYfshm
pxo5MWUrLqCcwyrc+bm5aaDOgTpc5b5jdHKWIBINuIURR/R4kByj/SEMLXyZo3D5
6G8mLjUKdSMIQAbUpoKDTNIYBAUA1S8rropL784e/mghKqVYrvokRYmbg753OXPN
czsQRA2InTiAxVqpE1lUBM7fr8FP1sfNthgBoefYK1FnnltnGnO9cR7iXKHLSLZO
j5Aenpl1eqmq/KbADH+yhDlzZqlKPs3HhyUsZ5MPw8b6IbDrSoH4P0+fkfRZxLGY
h0LTiQMd+C5X1sFxUTIRHg/cuwbGTRHXZbpxMLNc2kDNP8XBzd+0CkyCMTfCVW+z
wzyzWMb5k8sTATwd1xr/hTFrg4ZG9erXMiVLQ96beDFa6xFL31PyYqya2JkP+el1
2Xwm5As2ZQGfUzNtL/kyYn4j9RwSV0Z8aEK56FhTL0Q6rJi1QJyPpziCFWBC8EJo
bQLWG9Rz+KL6uyzeQRh0FPFCxrrEReXwsP50nPlwOhGXZ+XAx73t9HQLTTc1JEHT
ZqfeUI+fEeTJjzoBvJqhpqye0rRLTi2jSNtyWvqraY/vzCYE+FRDrTfX3BfWyhzV
VHfX53v9/c63eZ9CSWlQlGbbjxv73Iy3z0YM3Kn/iHh96ygpuMDEJiDM90lK4CoX
k2f02PDdcSPFV1vkdSCX42ydMS+DKvYZWHf5jwSih5q1FQHf79CH5sRYrrZbY7/l
Vyuu2JHlcgczeSEvccFTVdPeyn24oqwWv4Jlw34xRf211QajlPZtYyO5mYawY3+Y
iG4sKObnTZC2Yf1ETVOwY85++T1hLApIPV08ld56UO5K417WDYGffOxnjsewv6xf
edO72x+ftuOjJtgmTQok/CKjOoQ6C2aebNgkQRSAVfxtwvf1v9+s+3a0EEm3jl7/
zHFtZIyilvKFq3MFMz0wnZH29aNIO2BSjNCBfYQIac5uFYQ7YCn7P5mFbop11wer
3sdZ0A0IVtQcopNH5Ua3Z9Jm2jPJIZGhhzkdibGBwbN4XTIUIMH34p1whSDQGm6K
0fqAc2P1b2QKEfHojwX/CatXFux3ErkvsJSTAWz8BpNRjb3JMBBvyPysl0LzMTof
1RGMDmTj72/zZymwUkktPqTDgIGhHdo8vIg5cDsxdv/8V16wVYIHXUzrU0mzuUCD
HCKp0TrjCUI8/DUw3sXy3gKqr8776YIIGsS+cZK5hP9XfBNb+cO03LFTdPcCp/ob
HZVhJq8tmhxJxhn4q3O8IFjSzA6urfFL6H4uP2pFzedpjSkc4vF8StX30ZOE5/OJ
TvE4K6F3Vvp2PdwtT5Prat2idcNyKRNpsBwnX3Jkuwn1iqezZtrWuaQzs15c1ulT
k12QAiO6Jp2KsRo9mLoQzErR67aPIydDOIWWX9RMyGluvTr9UTvvrZiPQX8LYslS
1n0wysA/l8cp/raxfdHjRmSID7QVLDBTvHv9HPmcR7S4XInXNDQmnXMCQBL4NiHG
+fya4rzNtzHNyCiR4kbdho+6iBuwl1HYh0dd/U3rgTXAGGZAVfi20oDEv1Z+2qgP
gpLkyVBerWF+0OLI5CN1mqSuSrHghi0E/FrVt7ZYS3XHyivskFYXrJ5R/aYqU+Zi
4OkW1vFxUgL7Zj9kCepKzEgooMwdNHZfFnqyelz4EZBOlGverfxY0WH6jKgKoJGF
SWp7Gw3ohWOfBLoDPp/1tSaYJ2MPSpqtVQUB4ceVMwE/qhObVbaFoH7oDHSPNDXI
eMCletFr3lM5zX9dGwtXE/VYfsdDbKAdUYlGqZvT0dWzTKtCthFQpKruT8T9aLo6
yN6joTp2rKPtdjhzG0AKKLjn9bBJ+yZYT9Yts1hI9A2nJ3BWMd50H/1BJwsUXkCs
PYIjsX6TQ8DkKjkN6hqhRmx2EwYesnK+Pse+5znbnNBvqt/S6l6yz24FCKKI734L
BpImrW3dYbHf5KBLFZ6WwB5tGp+prvNWXlg9uDhyyws3cmz3ClcdbGrdep6UjiG5
YLuNSnYL7zhhkzgDaeD0YsRDqOWYjAS7xFk1FQVv3rbDRkMhcSuAZrikM92FZ8cM
7s2G+LmBGN8LQWetyl2LZyyT/o4Xp1M74ipEmXLWYHODzvs9WOt6IILnneYKD/tW
hwE9UVEZBl2PZgmctQcfPj/dwu0fJjFNyAekFizPG+xOrkXxCdrcI6upu95ELzRQ
BhFmk6VBYLDGwgb62HTGj6LK4KhkuUwemOc5CJeizp5tnJRz0ykwCoWLLPKNT96L
i0Fa1rQMyh/3aADPcTvJX3ZELp0k1hcYxdKuoSu8IT8SkN9i2Mz0B1LDZvT8E7O8
tPWCVlvrlXSgnhctgRvVO+7uioIezfwY6MBycWyk+6f12V2N/vAhSioELpSNlawe
WRx3ppknuW/x4ouyUxUkYqd8FbqwU06cVZtuHJjTxCyXe/wY/82LaYmyasKyWveM
bkTM4MWNYt3SqZH69JeU9I+R1S+I+aWGA1asNPety8c1VeJ0fDCB/HOpOlEG2AtG
/H9P9swJEEskuQsgofeRCW3+6g6lD49NwwGhCLreVUUfB8QzshzKOJaekM9jc4Qs
cc5pFt/ASeKn/UWowgPhoGI07lq7xxAq98o/0hF4oGWDq67ANSGGgLEmvknoIvYK
KAxL5pqR4urScqj2xBQ3e5gM2INpjMQSfmy794nlz2kSdju+8UGhMWIhGtwMGa4z
ciKlGBf2MbGt7qh4t5vrg6hnKuimbMNUh0gRb35WD2pCZJc35FaXjh9Iq7FJW0eb
Y3L8kU69n6e1L15CrIG3TamQzsDccpvt3LiudycpYkttUakv5PIOwfyu0ra/4MZP
gkc6B/ETS2aUgfd4VBjxkGwUMNFsVu5/+ToYGj8wpZxfNURrIbfcBZxmZLeqduPQ
QJi6I/QXhN46Vb9bUwXajkbINEOANyXTiIF+ZzzZ/0Y03ywbwhyZ9GRhxvQ8wRoC
DwsxzKihLrbk29CyAEDfKlMF/IRJj/YZTrG1D28k3gTltsmiHIFzQKk94RqRcxoA
rx05x5e2+DB1OmzrvazVX7w1U9rrDWKhzVRG+iPK2OFXxGujVodUd5p4luaszz9g
0B81sB4iCZ0CZuekPC1z27qzB4cZDzNEjTwdi/5zMT3QJIpmZQSDP/BfxwzXX8En
nYnQqjcU7TazJOau92DES226KMg8R/2DJCYlTrbBVpE5+eA7VnW7Ztq9nt5u7NZF
1JcSHAeF043C7iva/g1HRFu7/gtZg1CbKvTosJaBEL+ozER0aks/PKawwQQf0b6P
T4ES0UgRDE2Oce9BtduSKwsm5UZGAAHJVvJjKDawShayplvZS+lLdkixonOqRN/2
Otcj7SOoGBwwAHj6R6CeE8fLfUxLIGfkrC3GSXt2PspVfxpZOCi/9JjEslAWQptt
od12NBxXihJN7OCmR378GUkH4k7bc5P9YTDKk1Rnnyym0NZdALFFzx99Ty/lhJSU
XSVqwpvYS6TGj8cNuGb/evJNIgV+AKMMuVSB3QRE9170Fgh5TbbHgksVoEn4NjFt
GrwxHE/tETLaqS/DespeHJV4FukMQ9VXsVuA+6rVzFU+fc2/eZXh/2bc6IJE1d41
W4V9QZ/r/hCUnpvTC0yBjfmSVQb6UeWbkI0IM2Ul+8lR+M+7K9Wvev5stk+QUOOy
RQdK4gwai97NbdB7NlsaydOe/kLs0LNFB/wBiK+5m6RYYpkdN/40IpuYqINNXrCD
IzXlfNh+Wt9VmQtS1JqJKiKMUujxGH2/E17s4t3FnftsXi7A0Kw93lyBmL2YTCwu
Is7ULjcZq3SZQ87CmWrioE+yzVoG5uLD+ws2G4bypj0BzHgppW2aLDAoa2R0YrMf
adZY3dfJF49OjbXn2GmqMBWFKQIAEjONpW16XST0eBIQI+ap/PG6sSIRKOn9j8s0
D7ebqecPRD/hxLkKxHDDvZz06bP7tuPe7QGkn4ssOQZQTXql0fNo48VJv9q1EcW9
oPar7Qydxhz3pp4OfvA+zf6S/1lRiiB0WuM5JNcDdUsbqV8j7JajDMPlqIW8nxLu
xXREfZZbgDj19Sd/+kaa26KkW8orIbpTf58iUfXoUQt2vSw3GpaSOjRKQx1Hn6wD
9BSY9mpts/GmZJc4RYCPJ+VXDwBbaB8FOh4QhW+9+7w++lMpvB9ooGdRg+n5+1t4
GdCN6I2i9qa+hJsYMquR1LNANiRREaMFsABCeziIxa6rA8D/obED2mmuA9DxFEem
XmI4zN+HDh10w5TCU4esU8DQ5yJRNPNiL2OkYCGJ1/lx0qhkX3xdUBtnd//aPS7G
VpfpYCeXi/0b41NGIY+st0zK7VBJFv1v1lfYcS12LfkXG+x+74KEDi6aplkhkTRy
j8nVHy5dEi6qUnI7OWzlFUh8x9m6cqV3dGb7+kUeXyJ/ieemPPNLBwMm4fi9kCtf
8bvL9rxva70hRyoIvw3p4MV+Se7AI+gggfjIzHPf7i1nk+6qeqF8fTSbAztXUrkf
k+7lcVfsuaxxNDc3e0Xji657/fmVefAVLLGGbJb6VIgXFEAKHtZwrDu6bEEUvGme
c5rX/CbB2KVmSekc32KbtgOvDULMdIiJmdWIMYksgZtXHR3HNmPfkL+6/qPxKdfk
bXng03142soFA9DxKqhodGk+U5taTssCtQAmAKdWA2m46DjdtSOFYdQhn12t8vWs
7usVQfhX9jfkBKeLdH16j3WDJYtZLQK7gk9C8DagUuv2mz8KSfXNUnKzrobECSKt
C1moaEolLpjEGoVj76XJywRNuhMwS8WZWoNM/09mAzhkC9FgnWV22le6ebxKfXsO
dJdnP4TaZGMeH2A1fKFdLiluSW2Vg3J5A6V6NRfTzCwx/hdkG11NpIH1d6VE7gL8
sDBZKwJt5Po/TobUlxZNGlvZF0X94X1N6KrSG3xH7BVTD2GuXWay2YtNBhfKBFHQ
LBuB5+PG9x6R4MQxQFupHdZg9EPxCH3Zn5BPCFHdQbormahomT8roQ/VBplWI7Mt
05L6xeOmj5CvOLGTKPMZ+vLih38zaZA9AlE+dGxAMn0D2ScZGpW6a0tVhFAivW/w
oor40+CUuQu6U6c3HZrWshR29TETjSxFEIgQWj7z3dm7SMZcDRjXBjGv+XxBDjA8
rqvkQxomyQ2+Xt4/UCaK3mthydtrdj1Imn4sMT23emlGDLM/rqp+1ffpU7mXBK4Y
QODM46cfKgzlY3tamuoan8XI70A0PwXM9ajlcD9CjqC42s/2oBK1+XuyD9hQ7qG2
EpHx+HRVj8jrGjQeV8W4q6hqA1hL2rfktLQw+LrerjcVguEL20oW6R8SRY9jmMsk
Xrh2nAN6CRsTZESek740qOe/1ic6Em7fmop2ben/EEdPLD7YSaJlIyACgCXitxkZ
6qRY8aFKfNxrd8Yh/7NcjKTwFues7p6uPVkBeig7kvUlqYFLwJ9JLkzavMy8/+iL
x+QiiitrkiNdeSTD3k9uh86rxIlHlqHR38jWbPQ/n4W/MCqjFo6UjdVk4hWb5hXc
JS3trzQY6kCqtcfAiZ6G/wCOPWRpTmXcyVvA5hlzctMN6mFKm8Vxn2LMYyqDFvsW
HbktJp4250KabvISIqqcgoVGRM2eO+1zQIIo61LLcSFHD+BXuanYtM4ytLmm4Q6F
zaTmVQDLuGD9GSnzHIFGqIxp7CmbJ6U7ERk4Y8MQWIbDPSu1P3sMKTjr2DTzBK4p
XQA9lTB85kmlTnx0ZVKW0ztSDMNOZgpMcRbhddJSzmUpHdX1MdUXta5UyFHQl0D8
/t8dluOtRnvzh8Ejygz8qBDWP5l6sKTNKUuS4pWGNohS+9e/eZ9MzEjKlYJmX5mx
aqtKGwkQoyZH5IA2yOwN443vcv+li6R8LoWpWxMB6FPBzZTgKrizopeSytlSqEjj
OUpmpuVDPgiTHOEkXp55TVK5PN+Mx3+OdRHvW3Go1oaoafGUtJ+If/jdf6DGROH8
X8QJzYzbsqck1qpLvm4VGatqgkljM0P46ElFcfHfOtItn75Yb0qHSOHGbq8NuHAc
rp0bj1ly0JRhfaOhN1y9ONBPF/IbwPf7KBCXsq6LRU6dWmchTnlgP6ZG60DNI1UF
7TK/60JlLdy2JqqCGz7LB8QNq3JhWSWezJrJV5LaJIEE0XjIs4LfUfnX5aZU4InI
SKOImYsrshS8N1yu1FGB6iufjgrXft44/LuzqvQJSaqndJIj8a+94EfedwunA7UT
g5yns+iGtJ4Fh6SpLJRM7OgOMIiXr4uhtGhsZtFVm/UuqA4PNwl4PjmMdXaTb8NK
9w7YwGIyJHfVaIyOKdC6SLsfyTcl14bqQntVAoAlmRKv5OIyBCW0xc+yc4k+nMAH
NSFP18yn8svcnEhU3DFJ0uWmOGoNTj79K6L0VewKa2B0PEYsMsDfi3/ZkpCNZCC8
J10so9BDNnyPPKXUaJICUkTE+hs+2qSA941EUqhRYU+MZ5FLAGAhjCztFZAREAOb
qpjaBvzdXSxvtL6xME7bHJvuyBb9LDhdkEtosIgE/FgEGpZcFiitL5U8bRMozkXH
lYpPE3oYULkFv4Xpg92N3BEocGvPcC5CJFvPLhZ4WtO9F++XVqPuLXjKjqCXgM+F
kWALGS8G/Cy/LHrCjR2CkpKcYPp0sg9HjXIsmJHQdqXtt4lIPxz8w64t+XvOas35
QZbT5EJFUBHdM9m5+0LQwwc7azrKqWuJviTeIUM7Ps1mfp+YWDU8XzspoOqSppTD
M7PE+52p4+3CG+kQNz0MmPwAqP4eyDzHlDBbEJuBFh5RSrFrXF3AXxdSEtT/NnRc
Mlh+XvMosUjflHElRAQeU5JJ3dqWSWbbapgr7V+K49ls5cnFDRsOuEquI8KN/2u0
N9Uv85n3GRdwz+lIcQq/gxTtIm81IIC8pR9jS7b+3gI5K/lLw6ofGHqqNapGIH3d
HWsnu+3T+IJXGSymqYV0KxoIQXrHLUk52VSRYJkNetQ8zZc/rhnMRN5miavKC7CW
5AM2hQuAVspk1eU86JShKVdtad4SGWE8VLJoTFlmLQ5vMfQ545vFj9njdUK+6mQ3
xUCD+fwaF3Vufk2ItS1QQfa6CUiZOkdxcLP+wizpFlffaz4hAEvrp4EG7AjcNlKA
51CgFO+4oo+WIBJX7B3WObqADtSF+ukjqtXoX457SPrE07eovZSv6Ef4dF1907pA
DYiZhoZZ9xOb5HEWgQHQRFfVDYD5qNLynuK1GVwcjJIXnWLjAWEv5N4pfKEF4hL0
lhafZaQe4t57JYTWYjYNHBBO+hh4HRVOMsSjLcoHmleBWleT9VjGi95XDwBgKFou
8Fm83Hh2aaMd05rRxfR9eNy66O8wVS/zCE08lfnpL+tgKnDcxNbpFSq9nt8Kn2kL
wj3utDJ7b0GaGPTp1oTLlPdFNU8XYJdYx+ckczqlPdWiLWkdyOHWPDFJD6Q5npHJ
sxFQxCzT+vrtW8P0I60/ygccjsNVU8IZc7ZqDH4i5HLRRnSFB1NQ7y/kDp1qFM1y
gaUacupKDzCT/4mlO3xRx8mB7or8rMCECmKwIOh+AmGJnur3WiTR3NQltFlau6rb
mNvI+vbjQnCra93Ngalh4r/hmL22fu1yWWRBt4+SZj9YbkAarVZWklVq5/uMUUOL
HEQUkco6PUL9gtfx3hirUQ==
`pragma protect end_protected
