`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tqkRjIQNhf6CMj8+UlzFizpIC5S5BZHzg5WZrsNikAFsPBjkO97k74LJE/55aQSQ
2l57Fq1ON2aVkVl+ZamZlM73k/JPw90RluKR7n6wquuvve7oQy0yH/f9TLTv+gpd
TpnyptT0fyZiKvS8G+gQvIT6X0gQkx41KHyDTkwuuac=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15984)
ZSO37UCoDJOKqJSdPDZDXKg7gRYoQOhMhdaxbZ5OIh8fqYA9YdSs3P4JdiaVJeSP
/e5NBlAUIoGU4gUPzQAP5mtVYu5C342256TNhLbqBzL+yor3kYN+5yVhA20T2l+X
mKOm79I1sGahSfVzC6bGKo3sRxLC9Pu8q0F0j7bsZhY3EFhW1QyGd07fNpvLhPY2
gVWVFqS4pbnwsm0wXH6wpIUCVjQazMNERP2p2CFQsj8tVPmVZ5X7MYgTvjOrNB+O
VgpmUWTDt5UsAzJzA8quJuABoQPhWp+Hxw4D5nygQETFLSh1X+jRWw+0JZgNOBfa
byGEgqfOVRYSzQwl6CUd+oAupt/o9Lia95kwkwskrvfDV7fIhYfEYYTESF/U0iPI
PHL8QO5Qnkvpqt7tgAfeQMz/lyB/nm0Y0p2kxX7NITvXGm4uoOU2h88+RfZZMPFT
dQyXZetn93UNejuBqXaikqCG6Z/bSIvxJ0jUhnGx4x73jnwpeHcHsevyGpgHGenD
u2/SlwWsbFG7FRxsiy/WXbh7rwT/JsH4J7rPHsmpHAu0VT1kj+YY7JjpkbzO4ZqA
ggXWqWZV1u+V2c7eu1ScdxFushIFSYxZvDWnPltIAY74w5mLaVxQjAzP/q2iEYn1
AixW9ZoXkPBM710+mZpM2JIYRP9dg73yDn04CmWiYoY9AStgoftKyNZhbAjw8UAV
VmG8JQ4OZjPD+WB4ee76lC9STy/6p/3HRCWw4t0F01ZvnVlAR70wvg/kNLXzYmqI
ZVC1lVXbqJmVpvbNvZPEOyfM4z1A6TaDQqkvobuFiEDtzmz6+TlGWrH7g71akGaE
mGLG3MIwHshJsaR/Kle53pe1373loZZCcG9nrsJgz0o77VSsJ6XCYWW89oDAlF+D
5yvH+NuiQn7gKcdVXhbccmUaIscOYdbbGDwspf9uGIy+n65cVyECK76m4yMTzcib
D2SjYMSb9NKVg77vnncxlE97CVxc9SiBbEnRzLAxH16sTvK/L7W0d8sln3NAN4dl
SKw34RtK3l698dnLSMUwXJtIhPISUTnNPLbV69U4gyLtHyh4/NzdaH8c1PxBVRiS
a7IbecNeW/+Hv44jfWUk/7O1r/INXJc+3jU1aT9dcrjVXUVpQsYjonGGhOjlWImb
iGw5BjZ+SPUBvis8zsswJAdh9i6i3jrp93OZAfCXcKAuPzEs97lvIPtdnTScTu95
gc6zE5fbSzE7q+PnoNadNkxu/DQ0Wp7M3JxAr0Ia/JIA/Uxfzsuu6Omi1vDntULN
ymsVLoF3tpTfnfQQZU3eEIGvPXpFADcwGDEcYbDXPmi5EKi7odsW0etBVE6ksCQr
VvPJAskKKTbgyvkS8GBkd1NdCb9FzpJ/fXiGoUuWD6DBKdf61NO4h/KBx38m/gcB
WLTjmPFmHVa7NlJ32LZVBJRE4RwpzIQAorMOtRi8SUC0/aMkT+nQE/wqF1XpVOa1
koBMPWnR02CpLbhhjYwIYB0DYKQovfL2fuK9MdmEJP5ARDm9dxKyEW3epe/WW6MN
ccFD8bcKT/PdKZ1F/aC9AmxBhG5NGM7pSNbopDspr+YpPo2IdrartOfpcgKmDykH
lyXFhw155JSRjA+z6Au9EsAJ0/+Y/u9yV0WPFnkrREKnkEL/jFAGw970idDAjdll
KCrQZEfqCq7bh9hlX3jRpbg1rFvP3ut6IjASjnCKLV2iuwTUROulTjPfuXIrqSYN
0wvoitLBfaODt3aa/WhnJ5OfyNxTRLoUm0O/rZm5zWllljtauSxqoZtrl/wn8mbl
aO03TYdI1ep10HVSD0JOgr0kU0BQhzEFHlI/0psr0E9avVyP2EAFSBWBIfiadnFV
IrJ2hIxxGejnnQRZq/cBUNC4P6Pm/WTlirrAHHdkrg1TMLmkMnqxwo/OlzYZTNlv
YYXk66bQ9onE/r3Kg85AkeAUP6re636oKpw7bM/OMoz/ar0NRALE6OSYWU9cv7BS
MS8mPhIRvIehab/nmINZKQQyZ4yoIkC2GSCHKzbIUlmKpiF3vOfTkLY9gDUtWO2/
naQSTpN5iSpV8i20fwuT7UpSIOclxR4tayMGCPri6QcxlPWk/OWgMm2fHxLaBgkH
o0Z+r8sQ/dvSYOM1+AETLWOiTP2bM9go7zvxLxXBlNmHqygtc4tVmxajXjq1wzSA
C1rrOLPj1/TKTg+eTpwT4v6tC1vRL5G5k3UwTNJ16+GE0XEuu34uJzZMYQL7TVVL
m6jgU1MvoFlaR6uQFxiXuHY/TL/SMZ1NZ2CySbNgCwZoq+yZmgXr3Nz5l9+hvtAm
eBw35rhfXYgw978k8O62TLjbMGZz6QvxmMyyFqWigv1Br18kb1NymYf/XvUPU0vn
uajhYah9L3zdUquuJxoUGRCgVWcP6Dtm9FYY0JvF5453oQwUGKejkOhkPeTBPprl
SdQa8sMhIq+dEawwcphmZlOty8jeQ72Ms5qDU3MDWuNMIat6Bgk4htGX5mlzsbQP
f8aF8/bYVeqFbEbN9C/1MM5qqBvmGJmwux8zIdV3L3rViho9vqgCU29nsHqUfMEz
akQ1w1vhhaydXPaU7T5/JQHzCMtswQZDN9AYMvkBNtB21m05xBn20B/3DBCbuc4T
LaSaRCMzl17ciBgrzOCUkez5uaMndRCiQoUx0NAp2Q1WcA3opHny82dXKxyjYuc7
cqm68H9+f/1VE3DjJRg4x53JtI6hoWqwmVkMRe6hyK496WcpiGhdYH6FFqIY3b+T
w6KsMKwzy4UeNrG9cxeBUtP44FXzRbFF5iIRY0f0ONpZxWAx0baIYXp6beACYjv/
vL2V6IHepkrsVq/K9xUM7PioqGSwE2VjNjgcn+JZzi3LCYkQdzI0CrsRTvwqeqkR
xYarFxcuMfYzKVPH6m2EzzY9UIEbYsn6S6+6PPRTF1S62xUiESTQ3TPBouw1hud5
GXVHAKu8tSPMXqLHD2VCA9veWPTyne/Sw9N80dBefsfjHa6RxCZSrJMR0rjXe7s8
hzRnBGq+meY9U1sppvjorhpjbTbtQtY2CZpaLCHLG6gU9y49sSxSGmVn8aY/s1LU
CSdMlmT9yRK8gHReN1Gwgof0uh2Prquu+I8dlwQ4sceO7ixJMV0MEO/AscyXyvS+
INms34anDzh335MfBx8n7crXi/9g1Fbp+sNX2lQFyQrDkM6ZIWbAuWKzB6X9FKgY
gwQLmYX7A0/y3Bfo+U6liOSFqWtYngfWYk8GzTV6z+ctZUtu9nwFDTSmt/ZNRbLb
AvpNmTJc5rQIdRkuY6BfyfEsQ7/EHekbDFA0hnqWFWtCoctatt0vTaDWM2WAjMT8
kMwTGDj4mpxTmTKjFUUpmdeSn4YaFqAtsChfHTCse7wb3d+u85UD/wk92vkGEq4F
EFmfzSMjL5u3EH0JExkuRzKp3odHGYgY87RmC3LLqfzuLUJ0n7XEHUFHkh4RWQZh
AAYmAppB4gOJsw+PhMSUx0t4MNZRIAKD8pgUU6PKgtPL73CGE73NXtqv3awwSlLR
SxCWExWnQt8urGYfNI2ss+9KIPylDvI3siHsxvZWF4ctKw3yYVf5TG98Iw6jMvFL
krRwOHmpl6aq4AV2/Gu5+dlPLpad7efH1O//7zfNuEv4WUuZgz4LP9BzOglKrpHs
lblwan8LvpEMaySC7j6Irl7DgjHaNPzj1dkanzrg0qEdcwpvJx5e7aVC/i6dHojb
xxBYYv1ETeS7ooKNfUkCRNk2020SAbh3QR7mGJbKgZ6rNrjZRlbaSkSjLk7yKLe1
5zevU41imxQpbznjb6uv0HwZfXHOmbrL9Ttcdcecw+06B+05HEUpF389z8r5ZCJD
VGdtvm/XOvYULkRccITkgMXcvIrhSrvrNac5I0JeetNpuSy4LdG0c3fx3nM4lt61
dLyXob/YxPafHU7bWzMfi3qBq05LhVdTS0O8dS2ljvRc4Ho637rTwfr35v5wKzdY
0mHQHClJganpzhhne69KdGtJPxFc71fqLsjAHLBhvQ3j/zvEDirtH9XCwleIR9x/
4FkvH+b40nvl61b74isbf5Y6GqW0ncXrvtgGTA6w8IE2xRIpZK/25SwJ7+6jwFQd
wC4O+q6D3vbRmFIYDP1uHs1lryy2CHpDV2oByZicokQlbgD/yjaw/35V6hvSqjnq
4InTe3CipUyO7SrnhDEpBUZ00Wj05MYvMhGnJjNa5IIgoWCJM+aVrCOJ+dp2f4da
wzQZ1kF9ohDIWxdDTCdiVUXfmsLC/mje5On9kwA3+uOMxxs6tGliNqfClw16WxV6
wp+VvEoG7ungupq9CYqvbX46VNaA1ammqKCO6QWA+pLr+c1iFJBKdriD0SjTQ3yR
DvOuzNUrZllK4/g+X6Wu0lKFgvH27LbZryIV7YiC9L5Ngz5TnCbiVWOtYqIGXLYq
LJRTjxcdAK2bd7H8ZIKPRpAeEdJEdy5BbxjPykRuGwZ/risZMk3HVkhjXRM1IlXI
az3Cvi73aOosJ99Ux8EhDkcC3G3kNJ1koA4nG2xNSSjwRgmWA6/J9J97UotyO/kR
s2s56eDuC+xFQTkeTlXkMVhhGt4K8F1e99Pg03mlSOU0upVw1JFTQFFPi5mgZr4K
fOTuMViaOxpr3d8kuKAzuv29bRCLhnTJNtDhQt4TFsuNclP9RtPT5ByIx0vRKyip
QED64UQVPQvgi4itTmEaTJ3jekVChaWJyNyjT1IvPmWT2hG4yFnuxi3JjjKNsn6u
DNqmRR0F32MRQSBsJbC5yyWAutl3K7G/PzxMBMlz2Q8hK9L8uztVi5Q+SXhm4jtZ
rCx3489hANU4JOIHnSatbmANuAsmyltZGSFBmoACiz4Gve/fu3Yo17KQRP8zklYR
Ul6uczK0Jg0XVyKZEUnC/UItC2LYva3aotVrIIbPJeKBm7LLMLtRdgMTiAxDBsVL
n3szkVonZfFFvaD5C8V0osAu0RpNmR0RJvLQoo1y2umWSFCUeTdoDxGftHBN2jGx
fXEMXnbdOEt6IADU7MNQka/VCuv/qd+p2TNYcnf1STOi8PjtjYdXib+Bl/ISvw+G
Zh4cQ87DCmZenUZxu1/GocCZ7UDtc42S6esfWkMXgTRHGOWeYdGIUho9acPyQ3k7
4PZTRRxGVtMBWWTDIUavxuGzrltsixayNj7BiBLIXSmDqeRiUHolOkrvRBrTC7zw
b8hho1rViJ7hRJhMcPU7k8deMbwpuF2OzznKchbye6mQE4Mol+KdnS/PpF1mIR8V
NvDA0ozox/PqoseYTU/RUBnD1gLz/4lc5APmyk6ixOSSctqRsfNSm9DkiNsTKC0U
pR765wZ+ADJOTWx/ojmYQj0BVYiwv+F64QqRR56d/NLs0piL6BHsXV7hpJfm1MHG
AyPXsyBjUhmTe9hWpA0uPZf5gIFxhOyGEV1sg9fk82Xql9rBLD31N/YviIMsTw0r
a2+zKe3D7xZK2xmg8pEg7sCAMJfpWHmaDC9g1PLWCyflf4JeuskSO5IlDan+iUzS
BuSOzkaQ/n6HeXmlK+57Q/hkRmwGDF6snkzsE2GmUNkqHPvyxDOCStS0RE1AAC4y
KOuBNdJoNWXnbZwGsOcFhHCi62Z+HaUpTsJLIzytiH0+Fhm+d0AIZJkbcJ+Cl8ID
ZsrveWfSE5SSbnPipZ0r0U6p8FPUU1Z+dQ/Oe9RviRNJz+Fvt/ZW4n8daVK43YMC
0EfiSvPra/rmSU3hXQAGZw4XZjEp0fbLjR2xfpoimkRrX20+F22sAB+FRbrfWfcw
RaHK5zMfpzRWPWhORfxiTdItdF1sz/AdEmPSySlYkGNOEkyrpAtCRTnrfF8A/mFB
fjyINKqpNjK6K1gLbqsRvRgt/H0SxUlZM2Tj2sZGhZx+axdDj6VUnElFaxGw6QA4
ld5umgn/XNVSp5tYq9Kx/UVOYQj8XLnw63gurzCY/LP9WVWW5IX1JYDB4vzSmTzc
fgE4+744w8p1kh7jItiXBZNAgGhiIt6n0m6zWjsUFXXcQX+uVRsgIu/6HV7fYbmM
YTJ4GlDn+wszDNCax6THVjSzr3yPE+P41AuQMJpwwGWaXCOBiGvlztTVzU1MNRMx
Ta30O+uuMrnxlHCZZ+E3Fxvebv1lGCgMsEwyIWK7MxzPQz5QbWe3Z5SdX74JwpGm
1wpAzOfXoQjxMEqUSiCcOecgO2eGfFpRvAOMZ056mB4l8RYDvIGd3fLaZ5GHRMCe
NlWFw7O2eed7BaUjBxL3Nucl+oeMHd60MUzvH2JpxVk28iu1f098GCTX/JBQlUHw
rbRD3k4jUc8JVd/BYHSVxrL5YDC1qB/kBoFexrSwl0Gvuc0eM+tVGCxqut799ajR
9oynpAuCcFi0UFzq/HGJKGAw8bSMa6JDfNCwLZ7Ua26NWaxaFbuf9YahCkiX3JMw
hK1oE5Ri1yBeaFGrjvxc3/j5VmAh1KnMEaMhlhHjgcgtrIo6+SYVl/8JglEY7VnQ
9UwCId7IfrIiQuGrez6+MSbx2Iazmg3Ssm0BUgDGHcSMyR7LVAVAntRNpDvnWmYI
OFM6LTPRDzS4VyAy+vuXNrMCQ5m7MW7Zcwa3+5G6eQEyZAnUt6btFTwyraidTKY9
O+FloRIeAIO/R1DiMpYFZv+5W3OGDqQL8LO72kFtXaSHBOjuSftCQUcz/3NbWGWB
aU+CpHmcndHQs55vwv2+MZL4bVPKX1HXYCq4orEBBBUaSl39ihiv9It3XKNRNc7B
KnWJxLWPu2MbhXTQB6QPS/8xD4Rxb4+eFyz+Qt9NW3Gfljd/xgz7imAzu552r0aA
3jMDA6KLGuTS7KtYal8fZr+59u4gd3GLsQQkKyHizSQ1oQe0A9UJ05BvsEmPKRqz
b5DkQFqmSVzIeIIi0Isn5jgzN7InP2fTiW2XDNNnSgBhcKsnaI3tf5d/CFaStJg6
ffIpAL8/NK/VruoGeTreM2lhZTxjdIjw6doAi5jagSWL5gcLepS/Nq7gclWblmNU
Tf6GfZYJj//gKO335U79kzdvF469KZ+2AUmjXmQx64lPpyTpeCYAVcl3xDNN7v4K
gSyRxxUv1AtEefq/nhXFk8Hm23ODfjqPTSirshhsa8R2fLIfUNNk2112JWD8xMHw
OSdBnPr6FQPvaWNOHSKwM5gzyw+6pk8rf/uza3AObwDgR+bVf1vvZOPB7coSFX40
i5sLRiI4EyauR2J6CDTA9B+L+08otMPeqn1cVKzuLtFF4+IGH71fwTzU3QI5wFWp
KKH9VUlyhWYYwSVI3AcK24iQWsx+blBdw5uoRQNSW1z9C8Vcx98j92V3gSzYWB7e
ScseXiJuKaQV9l3OW8Aqkl/FiR/akPoB9+8+fDjMQfDt8jET6KQDWPKyMf6Enxl5
KCeTgi5ikRkF1p2smjROh0FONzA4232TCayHMmQafhVMUeFLiCrWNo19PXAZfg07
39fCy7PXVRdB3Yk4nJfe1wXjy8778lSi2LSDDD+qTRprxjzPDq4geBFo6iH/yTeo
lE0qTH6P4IGj8056626K2H60UxhZTdZ8JBfb/WT9k7pSkM5vXeN6Rd+OFPTRlAL0
U9ev570+qYalEezZB7kapAZ9QNQjPA7WD+CWVeW9O07KADQswrz8OsrgzZn1oMEA
p2mnmDZmWyvfb/OXBk/Y9DXkr9o/lcwZQso6xVXpTuVl81L/MR7YIlp9U7vvJqx9
iUbrJSdwyA6kCgcGIvBFmZ2NIUO9Eo3f9VrdDdwudI9zEF+Kb83VXOxHdNaEGATX
3j1ve8N5wS1M+HnZB8QXkch6Of0TnLEMW3Anrsdb3RWbq0HRgAb7bt6Sw3ceyxEd
euJ+GPjsAkeFM8t1o9qbG1lJH94p49WjS45jhTFcpDwSrUe+djUIY/Bu63KRWPnV
YUrCl8DZ5zAiJ94Xeyz6k1X3wAJwUG7+EchAqB+mLDU9AUgZ3CL/ymMOwkhKF/GX
ssTXFLY3mHSOfMeynuwpNvsxcUBhH9tDM+lQBxLLva2yf+HGihDiiUYhGKKQFLH2
2O61tWWp6lXWFW9vof91HU/oplYkNdXZ1ejkciHti4ftEuAVPY/GSTt/FoywfS1A
ywchjBDFjN8H3QDkMRYhAfUOVu36rR8gFsxFhGjKSb3oFaD1kOfyhjqqXIZw2+Q/
/uEDDEW4ruLSV3f5fT3VnBeYEHQ7eyHmvGOprBnwmRbN9gilS9ZmxJE2kj+h7yj+
Jqs4mOYwFI1aCMKJQpZn1jSMuoNaNRfA8HSSugpAzED1JzrpF0yM94+jmF6Wx3cG
BUshGutwcwMiqMM2GUX8/kbVwIPgTZXR8cYoG6pmQkumaJGJaDtiEEpMk3FONUeU
n88tj5UfTuguUtumGEIdGNuAeHhvQuTBCtn+aFO4SXAKBjvg5eb3h5TQde4OZGdQ
yUZS0H5KcVoNnemHRlhaVS+aN65XPsSbx+fiZsSfQswhcstUXL6AGEo6SO3uynvq
oRm+3ffCJY5NDyy1nzRHg6qZBq+x/qnBIzTNmFNdRGAvi3kMBf2LVgFipQlcI0jA
UXggryl6iDg5xi0aqK1lnxL+wExLnuU+rEfbLrhCf15UY+bwm0mALEVDpv5xeFDN
B9n3sgzbV4qXbcI19g5WV5aNRrrmoXy9/GfRkV43pu8ss1roImL7tlqktfl2J2LP
0HxAa6bup9AumRdDYsZs+Z7wmb5k7CCwg8QgkNDSKh4UIKoKis3EMFIEPTnVHThU
gC4OH4sq7zF3OmzsGdedGtrvZmu/MawuENjJsfg0SCTyPgVhojH+gkBJFj4cXps+
gGUFmZYqy+zQAvNz+kPAejw1KaH7BvGrPiuZ6YZ/+9LHezVv4Qix8wN0Kwp17fm0
LuB6LKAtejg0Rt1kkB0QsePYcY9iZHzaMMweGtfTsxSQ1jXprPMBzARQnVGtymA6
urRBt3eHZ6dXtnDm0Tm4HLTggrc7Br27O2fKrNF1UARokb+tv+60RPF0B4YUYlNt
+LqOoE99lFYMiD7HhmJQxqVFB5jvK+A79lzEshK86kf8R9puAinKppSusnHIsEKW
Sq5pga7kfWoCaHxdcloKIy0AUgkvedHqw8eU2IZDcQMXjjc0zQXEXUZoK/ZUeUFt
nLCHgVneeHJUpjfxYwSrgKbZ9t9Ykqv/BhqiHAzSREK7GFxj7DIDPx3nGwMGzkr4
XJQNPv+2K5xjl35LVKTbFO84fJLQlBEjdKSJ8B6U0ebPvKDIK2Fg4XUAlieGdc6k
NksWkS72d1eZhcB9N1uxIqTQuPjegixJ2t6+3eNXPDT311P2ZQgBh4gSt1lmTyme
LE6Btw0VLkbdDdchSvNx7ZShmZMdmMtNMiWYmZJF7Atl0AEsZmAXbSVIgphp7RDU
h4uQYvP75UQQeEnjqel3h4axI93M3UWdDV6bqHyBre8BcCgGyvQSMAhFqejKa9hF
dK8bI2s/vBvs3crNn+ed8g2oLx8SvB5ODBfoSwQuvdhxaBmPMaIzpJyWnf9fk/lF
SVz0WUAw5asqRApWgKteKDV7OEjv6I8rJwhBPfh8+aq6zPCAQ/d3zFggu2oZSIG0
yFPMuF8HnZgvPYsTVHZc2S5Rsk9KPSWiRsHDJ6Uc7hb/exBnBgJoeXRUc4/VzIde
ZDDnJfnyyksqMLCHoDnyH3C1Mj2YJUDDa1YICnvbGEldHqMFQonjKY8OvcpMBVcj
bwYjwYW5Hqb8cFRMT7pY2nAiQmakXtx1NhGcEaoK1iOqvfTYj/WiFGgbA+9GJJb6
XpBMqpfqieFywTcgvI6tY55lLHV5CApCtF5SapX0EZ/Xp4n0hlDrwpGkKjJdtkRq
jhtQOTYdYA16x0gCCWIWuGcDL074/yLrPwNxRSJmOYQU7cWS1SwpB0CN1W+TLbE3
3E9em6kcru17JiqLw/mfkqPQZD383IZ97kUdlmQaEa8XPognNyeSk1yszwvyj5C9
mvki6as7XQdco4Jai8tS0y8amu9mY0PrttF04BRRXZ+MLaQsuGRzqc/kanF5BreF
MpCaFtq+3qhx8jzutJeNkS39teAQuVmao3qvccf5oYdZJthLRzF1TDPDlxMzrrP6
CV/Rh2fNt5pYG4egrDlvvGcYJn61EpuP53+qz5expw9/VFajnrZY5LZDXI3LMUAc
UHWUJkFiOAr6hwh8lB1CSApoO3qwH+jn+4lTXoNhtIMcG4YIfOxuDqrA4avuAVGa
gMn/Q6rvbRK/2r9sWL8uKwJUS6Z172eXZE6LiM+jMRgm6bg5gSxm7Uv56KTmND4v
ULmeG0qydd2IdLZJWfe0yOjXNAbtFxfUI8Na95ZlBdp8JDwpMJx6BlQph9+U2dO0
S5OKJLmnpmaRo+i3VFiOB0b4NDu1PXI7bxt2QR1O3iaJS9myj3nzMiYGpFoJGGH8
+GtI/rx7uUiUicMBAr4PcvLDmZZy/HMfEEtJKjo+5/+W5p7aaIECl7mSE1QhC3y4
CD6ZDBeiA8bIGhDSyuxkJJeeAS1JYJa+gvM4ARuTcb/B5T+nJg0fdKqHLo1vHV6e
gAAolS6Thxsp+AOEk3A6++QELVi24aRGv9TqRcJGPj0XSfJA0Ku2FWJT6du1WtDT
fE4VFmDCDV2AzU0awmaTgh6+Qxn63Gc6wN5CliHDZmlj958zreazGddakXhz5jB5
+ivFcxOjS0bgD40fqpahWaxrvuwM6gnMM8CT9vEOE91o8LmpJzNkKXxYHzW0gvKo
I80Oh5fG/7663WIap2GdvFrtSkwJZZynu3aVfdlpeihGaKvx/Fd5bNElunNijpVg
miBt52ITpVseXuT64WFD+pFaAc47WzeRagHaSLBQhwgFtV63V30NYuNlits7W92H
0HMuhW1CdlIWci1MrYcKwCH5q7QLVoKOwRv1LcnLD2lyZng6xZI8qaPqbukyM5M7
8FAqi04Ee3hUbEem1SXZtssFvsJPBSMLIaygx6A9g3U1ZHdqlX2LqdYw7FD2Nrtd
/mewIZ7+TZZuiTcsWD68+I978L1j6MOix6rk6VW952y1Ws90qBF24yom0O20Pafx
sfQpGrY/nlHi/XpEtu7kwDBxnaYb1K3HzLTlISFWa/4TN3Xb9mZU7R9hlnue4JNg
8xp9Ku0vaKuQ2g5+SY/rBSVS1SZRg9b4sMhuql4ofQzix6OM5/+r6NzsWwcmjk/Z
Ct/myPG8kf+8vMbalOEb1/wU3Yl5xh2vvLaPh++fBwEBJJAGAxKjAM/yrlIP8FKz
znihsRyJERHMUeKvS2+6ZnQZ+EIWAJEdp4g772tw1gFIdP+lKnZwC70uYbqNxUXN
WDtAL7Sk6lVwBCHOzaRYq/ZqvBHqq9PBOdj+kQybyxBQDSG2nJXJ1yipZg8XvpY0
fPka95kD/hIuG9jHM15YkSi/kRXRrEqeMu3NU35ooYW1WiqcZ1tMwbfWQTPsaC46
GUB8dJQYxsA3a39tfxdSsMNbzi3arS2Cx9LQrIbYz7Gv71W6JGE0yPBYBDxKyiC2
z8Bw0889ubIEi5HAY3ZejQgcMKcF6NteuY62bVWKyxHmlHlQkCaiuvlGC3rYnFgh
+jfEirM6/B54pxSY6jM0w/NxtSwc3bFYWRWyBRG71tcZxfTIoqlrbDEZ1lCtiUDv
eueOnNPo8nQrX1OUnnxy8+DBowdhp4eJ8mWnmG3lSu8oBgItqXP21x/irXlFTx1J
wEywqsqObeGd8N7s/9Kdtvd1/2PK3Dd3Fa2AKYG27TSnI6vPqNKcI+8dYeZelwH1
8gAeze3VyK5mX72nNp4S1zOm++VuEZWKoKn6cqFXD232HGzLSEfZHXeTk4ztzWyg
i9q51VPkqrE4pQttfl2dTnNIN7WyLFrxdAQBGy6bQfTGssF4/ZfTQkKhg1s1vkQ0
YrpO92+0axaoGi9iMdQ9K0SB7IloBptR0xXZbNMyS+t2NwrOKyjwQTt8WBQgMAXs
pPuNEH7Gu56E/gK8tnpdy+SLcfsikk/QIW9CxbTiO0ZAWxn5rv2MNkwoxWMZmSH2
MWP6JYl0MoMDql94v6OxR/fiAGCPnIeC4t2mRDyhovPigtldv3Wo6tLhPT5NMIBI
ZKBNzn2uACKVBC0lnUFv9wniRf95EtjxIZimXMaJeDxwp/VVzzoIoV3MwQxWjMJ+
f1XNxLbsU2kMjZ2CPiwmU7VeYXscVywgcYUMnm0t1po1lqu8iHV8aSBLurGr5uxM
mOct82f6YAjSy1O/5OWA7ualsZj/qqMZiw6LUHZG2agmIhxQWedH5u1uZnVjJX56
UGojyugN0bIc/2909OiSZ2Eq/GNuTvPtAtKqWQ8GeMj7CpwlSm6qk/3xUlx96yo6
l0dxgOrbZX/iXTmBokcO+Kx6NyEC6MF0aNAypDEKbI2WfwWtgsGcFUg/MsyTxMXa
L50Zp5d90HY/89b7U/RO77PePz5yak9atdieiBHrg4gjfLexR3MzpPKFPv+msYfy
qlC8may4e92ohAB/PflmjWJyaaERdqpzkjHZZk1I1TLgqkmDpvMPMe8V/7jCgnem
L6fnUoWU3f49CjnB8cm3XZKoJjrz1MHTq5Tql3pLMu6EgO8rJw4brL5N3AcdtPM8
VbQbpQsHofkxNBc3mzWjcY/6f+OhZXDBez7/Zuob1nTb9TPqRXmvEKOCF/h7uifo
4PNWH2tVpvc9sVssOfEZ2+ur7laMfd1nLm/nlI039uzhp8tX/Ft0P/6yips8EbCJ
0VujWuM/Ws0LqTnFqFR0IVwNLHyNU9CbZrIvPg9EZqB/k4UHQrd7kS+CseS5uYrX
w4LFNWTrRJAA2fvGkX5MjxOvYoYo43iZeu9IbFm2LKV13wO6eRMEJ2eqzg3Oqjdv
CtskHKP1sHhTyq2q1iU30uIpmMgqTepNlqJFWN9mQTE6b7NqnKFtQa1RtBQefq/7
HqfBsN6gx/maIrtVJywFcB4/fWbNUKr5FUHYw0nrPiTSMNjrJmaAz3JqIHzVaFWb
fyf6oFO0Cu65P3nQZOdv2xBRA3sJcNlurhvsNtQCuQK6fKg4WD+ycqo5veSwngw0
yEUJ9Waq1U230xvOfAew+kcX1rlU9lNUttbCQm2qr4A614UrfE8ZuoFZ/EQHfbzh
wWOG7iU4qp1SI0pwEEs/1JhsEIamGqob2tZxnsnoS7Uof9VDskEVbBV4dEGcVz3T
/lvhW4fFK0jNvJ/D+6USQmDuwkqxllXzVCyOnsr9335NeKc1BW/AZ/+n+Puimetx
fjZ34Y+vUyyEtGzLa3pUT0kMYzPkm0fsGfCRDtcTvtqO8Gbs12WJwRTeA2j/9w3A
QNVWL7WSbkKQ8AyUHqVUBOzxjWdAjQ021+tmw5IT5ZNFj+NS1E4fd6GkChsstjNV
N+Tc0o1QMOQYa56MwdZNyuWNR2oNtQzWCFqfD2X3zN21FTrEdNaE2mx1FOjEKf0q
ztmCy9lsA1/O6XtG/1sKg0MvL9DHjP8WtPFtYI5PNy5RiPBTetoeqzCVcUFfXV8Y
kFo1SLxvMOtR08Wd2geVjUoL4J182p6zDJtXM7UHcHwOEafxAMnTBr01M7ByjdCf
5pv3Wt6spLB1d+trPoy5tqYw5v1y2olTXLWUpOkwHLvWUfV/WPorOO+crmYVSel3
cTAkjUHneWo6krWeiJ3lEpHcEWhBavso9iqIPCuxvnWasb8UAGO+/3pLdtbxpi71
OgmQExV3dPUFQ/oT02TX75aLUoz40W1YHa45zY/tmKiclzA5evX3h7NXfgXGp6AP
kEIJUcreAmzOFK8Dxv3gez3PR3q2HRddYKiNgab4BBqt6yMDL2GU13yM7fBJh6Lo
D0CG0tIfPvYuZyHyGtM13WnD0lHG54dr5mS3OYHI97pgZp4Awp4L7BVFFDCTNrIi
cfONQBLmXu575GhX6o0rkrYrxfu7hy/1LI28/SI1oT70cHEAhWJYDrERJX83YIzz
93FG1ZM4x7eKsGybMMNrBwOgR0yE1Q9w+I/Sn5MV4ZpSi+gAIojy+n8r9jOaEOwz
4xF2nmaoD1z+812tR4h+mhY50jdkUDFUhtnJrHv3rLKi3ZNVEQvNZXB68kdXTTVx
aKaiOCj4pW5I1eSmHZGVibM0oS0P1cHSFz9ljr9Td5VTwt0woiftS7lxr0omdF1z
ASTVtWYMlbq33oh4k5uvMLHvCsBipeKUHiTZvqOrc7Ub/cRmbPEXF1NwLoCsRkjf
6rc1SdMeHkNir5G8stpIV7NJBwRyXr0rYVcyf/ts5/WA7G2y03V8ouHr73nXXJmx
OjQvah4q2FIkI/fM5uwtETYfg3X/eXXAW3Z0zJMr+//Vm+6UMjTeriO3810QFo2n
3Vs/33mPeAviaQokjQrhtovFJg5Xgw9kt5aHO07Q64Tlcpvm2HrN4xKp6gm8W04s
myAUnDsAXggOa3QPrDtR7I5AeMKT0vxUp8Uq4u8+VKv2wghfnZ+JlgCG0XhmH5ti
rwOahlr2ddfY1w/EaNeUmYu4WEZJetGPGQnRpZG2MV1O7wPkCCQtmajRhgxuvNwZ
xVWkDVlCfop8hUbnjt8i2pzTh68ytqTIvHey25OtaC74Dw27C1EeSPnz2CEnh/4n
xPUhyYOszUAsHKNvyz4qpRILFpbzKvLM07JsgIiXo4onTNSW+t8QdbuG2uy6UJdX
xcsouvHZPilrTVpt9/lFetLbgjjVqdB4oYVbgYFglH1oPmaKTEWd1L8w1PWb1Rt5
ZtC/bL/3wrZHomoNSnYPLJCDJepfgpt3nBz0sJm9zeGcW7V/D73ZGHqkczKQbW3A
Pi75s/0Xd9mahXjRnv9OqgVnDqp9G2WkX0F5IzxSYaSkOD/fx1bK0nQC4yXYY9Va
fE9z3tWULa9isa2VGhJG4JKJ+6WgEg7qE+EI+8gDsSks1IhZUT6I3s3fiMYWLT9Y
58uTvxmh9ZnrI/yVgYMlBETiSKXA2jRKF2MuQLcWoYtAyH7ynuWXDC1H9iBqEJUK
kwv8NVwGQ/FGJ8ZzhEJaljnmLh2AqqOWv7VjkUDfE9rHVzZHWcokkCLnjmHdENiJ
M1ftLg+W71HclaKbhlHdXPgZTM0oDASlhwmEA7FcBeK5EUc1l5uSngeDUOUabqv1
UQKEcd5b9raF+uNUU/XixvTE9Bux56C8YkZSV+XRtYft3ghjggAXk+30tHv43oaM
sLwImQFFC7/HjaHhMqNX8Gr6GOaOjLJ8J51OVcUlNWmGxT17C3odJVjRu9F+KlSk
c28uSP7ifkcTF8g8X82u313hS6pfBcgrnvm6HbD5Ytu5lcothOJwmrrwslGx6AZ/
hOL7kPDJJwM/LchWD1zxV485xO2NiGQHfW8ehl8OikXNyhvg3utCFghEketzCf/i
+n/BCnMl3SLV+m7SYtaBC6BsMu1/2v/oecSAMMeoOtex/Old1bLcRClCPkXYfXuf
xYVTsoLRFXB7pBTTldUHbUe4fF2TBZktsVfewxkDhBBLYA9L8UQxpD/hrjAruP86
BWX6BHXtcYN4gwoTSgZDEuxO3OAeDrkst+Ys1Fz1JlYkaa9V7ZY+96l/juzISqQG
n9cz4thwqknI2ZEzWVEmPFQ6u7WAeWSF+t9Bo8Or26hM4y3avvC1Lttz0i++GwIO
uwY5tlIvNnyLN1SAzbIEtrBs67hoSaDTuB1jWb2X6TZwXqJQdUtAFerUEx+mCwOk
EsLQiiqKqJ6zrEoUOoxW4qyepJ6RLjIafkhtGB1pjI/cX6+SVHAtCSiLTfJGwfHJ
U5sGscbcRuXQdaHlNQD9ZYJvDvfdXO8avG7PRXWbtslpv1c0Mr54QFon/yQG5A45
D2IHOBO/IFnzyRPNB49q8deaOTSSmphpCUiF8fzUrMPUPaObZjmBn/qzZHTv4zWJ
RGT6XjpgLxpNyuOzF8zRsjLELWqXDLcTiAbpljkieAFEQbyAZF4I11btp5H///8j
P8EFWw/lcSiUP5kfaGwj/oCJAeiX0lff5Ya2dco7Sp6jrXkjzQruR0CTUT1owgwo
PDaBu9dslMY3R+T8jWRkrCNEodJiqLHeED/qpm3aqd/XUyUT4LD/1xaVn/3tkc+r
xBqv+VK3+gWZ2XuQr71pH5sBzx3ZgJfKMvEnZqulDZ7VLD54hqyd7asYs5SAKMK8
74BYTWcg1WmulMlKM4aJtN7MBD6kICDTCp1FuXw8SzTErusKePhjv5dc83GRiThZ
+EFb3s4t3ExtghMf4tWC2t76M64OtmwAvLBZW6UmGshE0sswHQbkwOkWORb3HIrM
a6TIB4NNNZtvrXSNkrAJbbDTFR5wtI6Bbsby/IM4nXJmUPqaogUzbNEHS1yUjXDH
Ygt61I1MdJWrFcySLEbBPv2QyvGZwcxyVTcicqxEBdmPe6OpTKH1Jdyt3/UIXWjL
AYtk3Pr548yzbkh8PHIiiVydHrHskI9g48AInSUsp4hsVhe2nPSzxGPBlZZ+qEcM
/wQ8hKn8MXdtxyZWNwGAMPMvPALp0H9sWJqHhuhSfuieJMAAp+NPNOPuJLSMO3d5
PbbnwIeOSqNsf+TJvBstTG69MkzNRqkO8Zv80po1DVssyJD/u34dMa5Xq7xq2cRG
pCZVjmXmchYvkkAwYzYJe5LE2mfgV2y3XOmJdEvrL0xtESI92CQwvHwEsDZK7v0j
OweP/bJz9ge6AWabJkZRGpmKHub+Mgogpx6Ga1J2aTZorWDyMnInYw6qI/JyYjJB
I90Hb589/uXRs7rPoJYjwk3AKK+t7xh0cQXan96blvb8J1JM9BfIMHdnWF0R3JtW
Moogqf9HxReV7Lum/qsnJxKpzvsqZ1ZynXnNJlCV6/19Y6Jv1B5NEraVcXPujlbe
e7KPvCD4pXZHPUkshu40je+efnhGkD/4CjtuDycmNEKNeISywrp1UOc/TT0JzK3E
wrwVQr+J7njjYtg9WTW5825YkVoB9prrFGD/Bk7JM0skSQaZeHqCsREha3l78caS
8vGslOWpBhQ7D1WhS/W4c31njH1Hj6UTE+wcXuTvHkmvZDa6TgPB938krOYbyXGO
rSM09oXbeU0FI3dgqfy5TbgZZGjE+z3idyFb3sGwUMymPs6bF77GbtSFl4TFmgf0
6V/LJUA/t3fPx9E0baBH4RFVb0n5g7tgGnzNVsgX1umHzf3ZJAiXXTJ0g1sEH5QS
NtVPZqeKxm+5GS0DD0nJKz2Ous7VThBXqETEKg5IdXNZJ9fKN3p5mYFtsLkBZJVI
Kb4WFViezRgibz9VnhLzit889YR4J5pBFOz2R5sqilqC8OfZ9vyoZWM0Ixz9/hWD
JPSOEXhDrkuaZaEO8q58Kpf0MsPDITZpnu2ic+8AtqZUdwtl9J33FUVwCK3NFPEe
DiIQNQ/Xwv/cMj9h+L2mfBz3jtY1j5NZALIsySd3dplMA+eqwVo+0oJylPZOHl+E
96EFOJmQIqC2K4grBHBzDYfiPHVxTSlDYBxXD9j8ECYje/uuDPGmJh3AiwUGM8Dt
qNDDqXx6wPS5mlsejIftCPVwPGXlSJAtR4uTmUrExBhY6llN83SPdz4vbgKQfHJ8
oHTJPyYOTGz4tO2kutf7jlJHxn5w5yKakS/nT2SYCmi+eX6TrVEZ/Xt0rTh8Fb7o
zAjsLWXYT7SszPXUJYcfOvgdA+Z5b5//7vTy4heQ5HNoSLroTT5T0UNI6tsASSq2
I9XE1MmAoVl34Abd3Od0jhBhIw9mSKkYit8xX/mYl0CDuOCvRkIf5Slv72NTu4kv
OK8Lplnp4YXfJLSMQccdeiVjaV17dwo7Ju6AKpBqaY8jZiCRvRstLjnYbpTBR1+t
qL/+4PSSOL2FHmtdbK4xp3+5tpBoN17IcCd1HGc1zNEEtjSCvdxpVss99T4BuJhp
zcYrB5ZhAr60RmxN16f7yhGvFOvFf3LCxxCQXTmDAipGhCIByNc4ynm5en8zObY9
gy0+4ZRfOmG+Slp8ofovPOI/RbOYIAdnYWJlQmtdQ+zRNbVT/kwCDa9ahKIDfcOy
yD9lY2wST2kpt62VvPAArWPnx83b5vYoOrmNUnHiZePOWKYtf4CXzGasc4UzMhJE
+Aj4rI7QJlE1rpJ8pMAueuEnJ1OZeptMEcQAYB/nzc1jkGYxcrfm6/xDqAC+HS0v
fJHN0kDPuNflsHEAYv0XuKRGFxUFGaX+mo9VeCPcuq7GY99+avrVypSGHcSTg8D7
zfcbHczxdaKtt1t1UPhzFKu6WA4j7iQIGjk7snZfnHsCLqLZVdGVErqBDAS6gdaG
j6emNuziPZAvbemnV8CkoUJyPPOaVflyISCuOecmb4EuKEIQ8fJslryP9ZKfXX9Y
brfU8slfnch4dA2EynwbBOMeEkRnRrr4dZ2Sd/1qxVZMURxZAKWrUGT2eXyv5k9o
9Hp/UTvhntAZnBTigh40eoZoDIgSZdMWu7samMqCmAQ4gd9xH0wGo4y5CNSc1m1S
MNry5H8HNpzhI8iIpsaod7b06/+1LtvbteKQshMS8ydWaP8xs0gl7Syx4ZpkOALj
JBs6pGi3n42cDaS29r2Nv6JLVI+kndU2RtfUxeMptFq3YPULj6SIP3KH/JETiR6O
U/Wp46kurA0erqoWRyBgYiI9/xL0F8iK2xuz6vi0XmLfBeCIOyskpxJGHjjnAfCA
VAtLTugpif35yJo/htVM/jAKdacj4p7bpJnAIlaXh2pqY4aZ+vgUCaB0JAkfxa/H
jRp/RxNbeKqmtxXG+f02PAJbMthc/lce0+RWY5k23u3PSGQMYyUfyVwDTOSRVYqC
o+AlXBzRRdGhgNQYsRY67orCoOgr+wb3H1d7oQS/NBK1Bpv7vf5GNPaKIqMWKFKZ
9JqqsC9AfNyma/gKPxAOyHPyn6QJIM6QkXXrKNaguHGAeaZXk/rACHaP5w+zzf58
I72z07TuK+gV3WiRz0HFSs+z+d5Glomm0os+juRsesEoKBYH3hQ+uvfR/kSsV2jy
bujjf2O30uR7HopAljfvREIJ275Vn7mDc2BE7cNA4/Qiwa3xKvdlMxHm36bBNO4O
j6lZOCYx27FWNhnDK8llRw/ZjGhRqOg3mtoAuRhQue8P/OhRvPiZzWPWDlXhNyRV
4S/eU3NvquZ3+xq+XOW/dB+6S9w5j1JdqymMGuGZmwyHNljL6ufAiWptxkcrC0hK
CVA3+XZH0rh+e2osZEVJ/8YmZN8zKNaN5O/3YDVn0+w3vQ5uzXREOUC9cD/ucHfk
z/qY9Ns2Mq05aTRdwDZzpyaYb1RD6eTk0d0VdyR2sp2NoQ+lNl1RXmmN0WFvElKf
f/bgCJ9Awy1m4dLdQWvjb7FGZwSbOEvAVaBwrMu6EgLp6pZFnhmGYzUR3ZfGoyEm
5VUFBqq5tjIuZJ/WX1ANuG5FEbo5hEiszPwiIc6l3UpeSl912sU9757QaKi+19f4
OkGC9+HzFm7gpQKoJHJ28g0Elonf71KIneEPHR+NFZcQMWTkWNQeDF4HceziGsuf
dijGuw0JFETpUXaGhLejyKRpOF/kThMKfoQY/lz6fYlY3ccXeUjsJeTedHd1K9JJ
gAQeGl55EhmxowaNeMpeZtGkFxsHbPzWkTGaxL06E857bOy5qWFn7iEiMjUiPCdK
BKF/GRruuagl/dWwR0Ng43rfsby0bWcseq9dkExfFGBZJFzqtI+aHEi/rmBkqUbo
BeY9e6KAaBdNXrGa21VR2IN9E+UFFmssgRl2ORLMMhEPjMzU07Y8PAha+0hhWr5R
kG9lZU0D+ULfwFVprW1vqabyGPPBeoTwfsXsHQjy3GZBBvaK9EJd0vgb4kt4hU7V
LNx7KhmJAQoX3TaAcSBzTuMVPVYKXEuhj7YpfBDSCsr75qH8m615Mg95qZezOsjs
tyiUk1/fu50OykDLtcUvuTUFe7nzUMipRhXamUqlDEZ3OP9GBg0bhgwJe1jh2N6N
MM9K/1ewSsQ5kyQ2WH8LEByKnlR394xVJ2QbNeTWwoDNpjq20X52Fos6fYaEI57z
iG5qtJMd1GcnHVD1TiNIIJw755SEhsImVJHwOcSrW073KNunb3L4HjSSCvmVNkUH
/OhBfbkEg7svakCqgMefwzMg4A1MaejKQ13y+4lF/umP/+JHa4bps0awgeH5uIoS
W2dyWpJqmr2Cj07buGMckhm49H0O3hA0TGTMNrUNx4NIwbVds6kgtOLpW5/e4Lu8
a02ObByRQiZzJWr2Lr1pg1RyuFAOlCDgRbpvLz9evZBEvkGmjZmzch39Vw7aLdYF
o62/D0/5zWNenMIhNly87OcVL9hXSb6jPvFLBbtzBaS31hHrfCdvuEzuYLuWVpve
/G1xTo1awdTrKYl2K6YjT/SVBny5Kqr5cj5SFHuMBuBHWp6lVve0/5duVRC1QlNJ
lWxMDduEYwUYjOETQgip1qVEbkuJdDZXrQpgITDxmx9lyg3nC7VuuIVkTDTTHiUv
fXeYbr4A+1urW8jYA9J2U0y+fEBtxXQc+U7iwOdWC0TUio20z9JsE5e2S6j4fPQM
TO8QNCxOZBcDViu7es+Kzgo8rqo8aGOh4aPKRkMwxsdF8e9EbB7DsSM06WPHQJ8U
dEFFnW1/gqP9pNsnxSTldVejNL4aPUkH4MoKs7hEq64TOzEwlVrLAYqSoL2nlOHz
UbKvPU1qqxYxkBegfia8PGCGJBDP5gO32JTnrCPfHyBp/p2ser41OqzFzmdayztV
bLGsEp0OBD2fJl3xxNjlBq68+gJp/slwPkaq2ee/qILWw4Lv2h5HFE6GgBUxUNU6
+6nXXfY2gCU2rHW22aMu6BZZvhD/SRpGqLR/MK5dHvz7bjOUKHeVuz1im+r7y9pY
Uv275qZVmYPXY4v2UZyadUViDc5JxScWKljioZhjOdtT92ebstTOX66qKrkXAXRT
TaoCtzqvJvNV4V2t/0KDwNl6r3ai/IAbsJsE7FO+h6JdSdfYG6Q3phoAjvpIi5Pb
tD/sg3ZJpeKdkJVPFWEK7YfaehJkTKqUfzjg6g3w5M/8WvJDDvZZDnumSK09PtlZ
vaoA6+FsviwzGcu9Sny5pG6Fb2SawfTcjfZyJ3158xk20TRDk4egZTzUfRQ6ouwE
jRnGhzMsuFZukVlZAa8AF0dsakyOFP5rnH5sHSKPX2hmAjTg/yWVsU2Q0SROsJ/P
4Cg0yLHInhN6e9GNAt+x8YB7aReHTYDA3abtjh0X/qw5IbO0O05eM9EAb/dn8k2r
WNUlD+MPFr3jR1uj3XsioW2jgAF5q+rBCrs/XFuxyRbW1KD5URsAzhx8cZ6Mm1QX
w/cfPO+lJHSvbw3Qc0AgvtJHbcBCuQuglzp80b+rr+MKUYU7GWQxGd/FwWOuiXb9
A3hIDpMvUiLOCyrje9k2QfH/04LDizNbDvZSNI28yP0C2e2NqVr/C2QAops/PUE5
`pragma protect end_protected
