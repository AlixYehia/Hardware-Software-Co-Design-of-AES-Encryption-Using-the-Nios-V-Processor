`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dt5SmhC1MY5Q3MRXJHVHZg6vQ3qBLBsvlaN2LQ/wiKrNLjaGBLIpkJJ3Z77NSzLV
1NPxwGEi68CspmLIW6Vw3NcGMQxAwAIw2PYY+vbudRTHSnAe42vYQRaEmGgywC3G
tQc8QHmVTseTmB7Wfwz9YePMdnR+k/TSaK32cSyBV9Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11264)
OwXzG2ucpGaZq33Hd2tSefRr7LgAUKQhesqjXoutsGiTNKiY5cgCN4EzJTyKX5l2
/fmUt8AxFRCdCSeztqKYy2iGkQVDI701+bYyXOxvJLfD8Iz2XhL7i/GhXXfa8sVv
/IagKa4xJAvpBS43VAy+WeFIUZTxT/gYWf80iiOyYZ3XVo/ibpytngcJg/JDbQeF
1uqQxD/86G/klpykqHAfifZ7Q4Mt4XPnzMpCyM1ucO4pJh/YotzeIxmkrWt5Wtbv
NHnfjDFL+dOwG2Hde/LhNXSFcyr/tl9kXrFBbkYplpePCBtbQCHKA/FCT0LUCcmC
0uw6ZP9K4r9XpSVI4tVukKWWXaRufAeMGwxckjupv+Rayyy5y4ZQg4pOpaA6Eg1n
lywMsk78LkH4ZEmPxoVelqX7hKebhPaF01JCKf3HnrHJZ6SzFK8e0+fzwUTlunxq
zla3k4kHK7ttFNvrFLU7GY7hfiMK7coiPrsZ4aYfg+bJ34a1JBYrscEAuSdlfq1C
6iyUxpmDBlkhhcSJzYlV7NnRi9lsFr0o5SZQrzuESnNoVk58nZ/EPvz7vMW7oZ6d
GZ8LG+C2QOIbDUMaojSk6rAJDSCLHOIskwUzL1ZUCR+ZyOpD+iNgdoUK1xMQDKCd
U9UAbKyfHW6MSVHwlwmBZlwfeII601IlXnRFjP//XSD4+B5riJRqwz6KAFBHbfu8
hfwX7Qsr7ItFCyeCXjJBMcKFaqKRi6NQpJFbDFZmqw35i+nTTCVX6CezodL0hFUi
lH4R7hy9RFM1oAjdI1IRRsUcJZzTRusU2EiHOV8P3BCDi87OwGjqGUbZjXovEieR
zvfmQYipoSMg5KaAZ0Dujt8HPRzeZryjNDJaNtIG6j+F5YK7WTG+TgXdEEr6ugfz
wmgM+UFsVT5eZi7UNPHoGgSo/mX+I1nDvMR9yipWB4KTXrmJg3gminmA039qJvOO
Zv1BBjwDReO139bQdFLdqFlunXwR3jwEyV8A3Cso8CeJDMLnkwdUq7it/+CMCjBy
cwPqXXHsN48k61f3MMmaI0LwboNYF/n89curAabs6OTva888oEqq63whFFMJV2n6
KxdinMgLg13SPQRnGNa3E8NqYN6fe3PSW0XUkpS6+P1txB7oW1xO3u0bb6txHDfa
TYc7ga2I/OSqaiH1JjFss+UDRn/hpDAxzUa9UKsKDTJnYKARSWj+o+KOF5ptmHfl
jCymnEQoeqUwD78srYPB74rQi5Sz4XGvLD1WW0oly4f7CGm3IgJeV9x3lr3EdgiM
CMAgOVzTsetUfZZ5e0I0ILOThfuEQMVUvGASVpA9nvu9Kcv5x7QwKAudEhg57ZoO
/FiwsE4OcjkAOWgBiuoSEih7jYzbnJKuNZ6Ss/l/PmPJa60ogs0WTytdNOOhcg+w
fy6C9pRWJv16Z9N+AmKTPDHc60qhT0j2XJQ39z4vM7Xfoho97Tqf3JSH4cirY/B8
pztmWXA5UAPwvDDdvZ+6YDMMHBlU3LRg6D+hvzy397fA+5nZzrs7VgTYOGXjZDln
EEfRQKSntiQnwTScx9QrQBA4EJSb2pRQtH/mOHX8Lzy84ueuooEvyVV4VlWxSyoj
yzZFeWSNA6VBy8BPqo9lJtO1YCX+sVWTbgbOwL0gv9/QOkUAfO960ThEo2fGnf/J
74teoTr+BMS6F/QT1OhvD2Z9/XDgR42L9gR/FGHTBF3jbbV94ulD7Jla5xgtEOMH
qk7sF+oWAx75eXbdOlQtDOpphJ4F4uN76jh3sNYEaYj/qqSLjqQZDKy51qZ2Zmmm
qFjybReZSq/rNV1BQSEmp/HSlB8W/++d7v2IBbMuJL1d2VfYwvAUAyMwZ7RhOqgT
0KJhZVWlaMK8/Q8gXTVqyC9sdnvGrvcL/AIvU7Ylg2XNXWlUUze53pVKVnI2h1sB
zkc0IN1ZSVAcFArhqUMNCso2qZ2NVqkCR2m0NnAVUgr5Ls2t4yxf/UaijXGN3Qhv
Pb0bcYuEhgxdpkXzuxeMZQrYIX78qvhpI2DGkgdeqDyxeYPHj67yr0SE8bNS8OC4
ccy0AkeUU52O10YrWpt1BM7PPGRWnHOWrd9eXafzKMhTnPLVkagY/Fg4l0cP/+n5
vi90mW4noeVux5/LFch9K+8Hc0AgvhZ7ixESof6t03Za8nxBPCUd+GGQ8tpSc+4k
xRHcuPXyQ2bmU+D6ng1OLVxMj2/KfXp2eUtNrtc9RUDVvp1Y9xMlutCUL/RwmsyL
kdmPiTYiJaeQbGRg2+mIs1mVt7j1N1RYjNM7XhalZXkfTCMT14aBeLiYpiYfM5bC
gZyDT/Q37FnGwVKouS1IeCsMOf3EfTBlP+LwpnN5u4JXbOZAcTisXInBDpx9u7lM
EIGyPM6h/h1h70uyE5WcO7rSGNqj8yROtxLAHS+DxSEeJCtQuH//Y7+0BAoolBTI
xeDxC7hcfXr27yLgpMLZxwDECOWyESHPqQ1JCOXTAOln3OhmWLNImkeg/ZEDXl5c
anDfTDH2GHm8DQprqoabW79wGTVu0FX/UUDLSZ3VaEwDrJQhI7nriv8MbxGOwE1b
FjMAc6guQBEugTagsd8xv+tCOiRcqdlI2RoTNViO+mvUpPFpIcns86sfw5XHfHA4
iUyPrgT1MM9woFFHwVpmR7lAlsIKHnnjlYfsHyGYvF2jgD8gngELaJH8vUY6Z3rS
d8GoSL84f1u4AmiZsI5KwZGgCBxPQAFhtz8nxVmb8MblWJZUwj+kdik7WE4HChPf
XZDCEwpPiza3jSg13TNaY3XwnlGy20wJLSlFD/We4GmgAFpcKV+m2iYGm8HJb4xJ
Ggx+myMLh9Eh60N2STMcCBsHfYvvklIrMj91U/TkUgup+ouj0BSaQ2FP3+TvBlOI
mtO1wT9niQsLJiaOPUP7ExhQnHh2tCAe6i3W0c1mNs7sRPOxW8pgSLpQUI9Kzhtq
K4SuSLUdv804IjmqzLakfZ7FlH65jy8zLPr6Ufwu9sfxdr7MIgIA7wbpxO2gYspo
woE+T6JRv6kvOQKYCoVdHW6W9Q6A0UHCW2ZzF0P5XOjLSSRvyG9yBWzs0CoUjr34
XQq58Uo32v5vDApD7iB+IwmThQMW2zxdunS5vvcxw8x+6lkaizjl9fiS9XtH+kNo
6dRw3uZ5ZU1yDo3+VFeThCqDBhNzXK1S+NQ+ADRJPeLAzZzVB4x2H300mrGUZpKd
+QKJCoSS0wlXit5NfKLbk2nscYYeOrcCk39DIvGVX7hdc1h0RAe2gfarEnRELdfp
gTBZ3cVkp7CaaM0jBUq3hbzZAMBblkJT7pyiqarnzLmZMFfUB6Gojt22VTqdeaim
gGzucBNenpJJYYiI67CHR2CzMNQedocqCroI0c26RT9KzANtPAYIW6EF80oODZS6
zTwdQOQBD88osiRZQmR4icI+fP5Hgp+b/63+szulAF9egFmUyrQvojV8Eb0s1s/g
+NuIw65RZiX08B5x5XhBbtrtKp8F5IFqbL+iRSXKMTMwV2Z/hpMNkMG5pbfIKuGA
4nx8Q5AOW/lOecLbG8SQt41vln9aB7H37k3ZDMm0Dn5t9D6c1PAQIsYamdwtljHk
didannwzMqHVaf6hxLf5081XNmK4NTPqev8d6KanOVWBwV54RguiwFWKhRadHErp
Qx42TRSiVTORaH5DNi68BAkWZc0H7/5k5DVhWuc9OjYNwn0cTPzJdehtYTNKk0U1
bwP4TWfrsPFbKhvf4+/uVTBIQIuLZHP2q4Y35cs6/3fxfI7TzUuUTKYwLPeT1qDL
UzR0VMsw1zLiLTDni6ZTEXZB/4P5GzJzTRIuQj9U19AS1EnBrqUA2UhuhRlQzGIY
OQQktLth7RZ+jdzHYNwYbjuE2ETxL4h8PN1Uj4Hc82nuBtgWsi9pSuS4KqztGDwM
oaNQwJY46Fwv2QQWIDGQK1kWQX+Mqycwo/qlMUbTXO/hbAiLy71agpT99rWyitEF
IaiNMZqwdauYIZGucZzRaEx7OAi06euUBUc3XTEDDv+8mrUCPMFSfFT3NfPzh6C9
DwCPMMqPNG38DEPbqOUJvaS/iAl1cP4c/VDbB3I7bZ/jb/Fsgz1oR1ZAyINoL1kw
Oxs2JupjD1/ocMrEUNAKpyNhEvg0KS95M91jMNVDb55YVmbLNluBPnuagSktpQLf
cSVxi4jO8OD5QqiTS+7qBrlPCCSbGF08ilrRlIMDdUh3/I5kJ3iKCNCU7SVa69xS
JFzvQ3tu5/or36c8ZfW+2LR1qb4jTPHxcPHJDEfaAwz21z/PQrAIbHq29ohv2Hso
LfNqQHnuEJ0yrmbRhsg/r0t1JYYzfQTnP7ntGobuzgFsWINd+myjcn80SQXmAWu+
bCyoDHS1A3Og3qnWdWLzqFNTogNWaiIOYXmcQWhAadSa8KxnaO0oKz8bSYLMMDTD
GhCEkg5gTE3lu6p2KjYfY4+TP3v15TmeUzTrWg+XHbBxOeXi7pt00DX7qel/PL8a
75D4SGEbxJaSwEVTPzyMEJgWZoW70K86+O/NHxuCoux4Ts0Jto1qdMXmq+tshqAa
WKa8ICqoediA+e1Lu2PV0Qm/PyDsk/6TdqLiujNPf2LTeRX+BVHxqArnSjYKN/5V
kTFzgRTSN1EF+9q9Blu8EtP51wKOyKtUKvbKb4W7kq4jqLbQkhnpbQBqlIhKmbvt
G9E3gefRSedxABqpu/SmZ1gxbtO6SxVq7qbpskgLqCkcDtOfgiuc2oO4S7kuMCpM
n5+Cfw/oP5P42pZYpDBGxYbvUGBu71CgZzMQURHMMFSr9B5f22lNxk/erHpFVc66
JeQRBbtypIcx0pFpizHo4lVyDQniSFKPDAeVamOK1TMnXAbWoHvAEwCZdOwvuFqw
yaDSiYQ2CiWMA9CDgqv6/Dbgmt0RTw85RUliQkMbscoVmnx5Bkug3YHZIi2h0fZx
lamCGMn0rMZoHHkKmt4TY9qpWjrUbv+hnJt//7HSP3TGB9jdq+0WBalk/nVd0I5j
bKxNeKk1npTW/ve5jpj8nzpUz4z2tWpTMAWy0WI45fYOvdFUrmNo4ePTIgPf574v
GSYYBPjwb+41fcXcxyJkgT8Sw8njJ87bavZKMNsLNS+mhw9uFWvN0VydGzY/2A8q
weuW5ydzIbQA/hkShR3mMX0PhzkITS3/SS8Mp1esFyVeNFHl0xmoggCsWTLS4bPU
3czU3ZromoXtl5j7gXggGGG8YJPgEDlGC6rJZtxn04eksxybU5IDAwgCtwyfoAye
oW1BDBEL5K5PacNAlOG+wvMoBMAF/UJigqYq2Y8uy1kHorRxBMmfTAbPECYS7Xlw
nfLj7w36D8aVADiTiV27qRADxM40yhf6kEX60gPxku47CX9nDbjKd6M5d5JBf+P9
j8rPcDEQHGbcQP2UXd/1vHEclgQg4/BAxNDcrzRUFLNMfSuU+VBgdsHnYCwixdS+
VbHciEYFfac2mJcMXKI/76k+wnNNEKeQTjZ/flo/0NPrmULXruFwAnz9HAzwgfe4
KMJGIfutfwwH9LenfUJoRWJtQ5n5HWoQRSOSuT/QJjW/yHkgpebDv4AeCZQt3Z5s
F1SI8PYNFEi6j9L8bmsjMe5As3jgIgZ2C1gO+KwtzV5o1WWk9xNL/UGTAccy3NfA
nwQMpHcmYjyYgqdaBx9mLSgWs+Wwm1D+BkEnvzi1i/xsA5sSDsjYj4u0DNsA/3dT
4uVzQe1eY1IVFV0jrxOoqs2rE7yP1GOM1r4CpFJnY+4KlSgEuw9i6XwuilZYiGdf
+l7R5AThq5tk2fwOARy1qN0jKC4jqLwBUg9AIpITh57jOYErZ4MSfVwk/JOCKPg9
0TtA2mm3jucLEli+PhMvWrMuwCPWPLsNzSOShNP6G1HC2Bqbwg1otJDzVXC2lvel
CeTCLTbJ/9YX4Ww6YzhZDHb//btcLG6Trk3b6fnUhAQt0zE8Ob+axGQvLLygifIY
dPB3WRE5QGJgbxrqJ5858KXXoM/GABmUEp2+JfQwD3wqPL8PcawLPfeVxmmGi4ag
9NvdrifhnW2oi7c/IdAhKF93HwKeeMHASo2LKwlLkpTWPPcm2sF2nt8+dbCgYvUU
oCI5FF8zhJwldSFnFob+5ah5IaUuqfmHeBHrtVG/z/IrUV0c7DQ2yTwJCayii3Dz
ble2l91SP6H3dSkslKwpUt+fvzMBAxefQnSKMOqMoYS25Yc8MjxmrMdje0544E2G
FpmmMBBCcFUuzfkdkkezSj8rfZsFfIQykrQ8TLoP+ojw3pSf1dq0aqDYa/BipYBA
+UJCFAPFQs2hPV5PBGj0BgTd7/9CE/fPobKb2XTEQmK0PrYUwYETjns71sorHDxo
51gxi6h5NUX9yT/RlAcgD5nMRAFtPB7DRORtEIuu2qOrNmIXOwcO8DBF8vwytfDQ
7nJRBBqCXj3eezK4dyb+2PU59dl18qgSIrsCEnAnKTRJXH6hFxbsUZmsyxy9uVwe
QrvxFbQbulTM8VXyLv7P0mYL/s7Qk0R+6MsOpBFuDT1COtnorgZmJxpqjZbZdRMW
qvG5XlrAoz9bQVUVc5ygA64pmgxGe6IXgtP2EBcFACLqyaSup6uoIONvLZrQW5YK
uUiKGVnizOF2ZVN5LVgR6tJ1PyXkR2NvJfICUMXgURdNxQ/OeapAciuvB4ipzIgH
t7+cpZbP2R9JSPzSdWks5yO206aP7SKMPrGDvfG2Ykade8GQ8QiXpoctoIyGlllg
GopGGv2Dk8TZIA7l4iEXCSUTwaDrg7ksnEYW8ux5R8LqSF15lNs/zzy83a+IfEL8
hIzK14Wxqg5q3U1jP/ssnpQX1G2nZP5iMh9VeKX0dbeEG8ClkvXxgIC6d6DONT66
xnknd7Mq8DW2V3dzUseezugC/h2uNU12pPveYh2yfB5B7QIQ4TyiEHQISAbefxJt
VMM0hFbZj+T/Uz77qXTK3AGfMQ67rC6Zhv7z5Pu7aTUQ7NZ2SZulJfz0tV8Z5lff
W62X+Za51/hB4Dwh5x2udZG7qlQo0oxUWiLrLGJwC1Wl1/HIwDqUTsdO5zv52FHt
AnSsY2NPv4qvUHOJV/VIAgNyWgoJPUVsddACA2I+/WPhprRe/fzc0+2C0JqqxaTU
HcVeVFZEs6xnm5H570JScj9DBmgoRcexAO7+f4qC0TDv5KW7FhLxlG8Rem1LRlkq
yMe+Qd7LcDZNjVyeYADL6L3beTC4n9CsqtXdb2sAjrJi7mJtZz5EnhCi0D99J6Rq
VEkQS4s7OYi72KnPUBaJUzzCcXQv/8/tiGHAMGl12HhK5UiBwgoA+bdPeYtmmJZZ
4FXgZ4OL3mv4PjXl7cySN3s0ExSUEd9fnbuj09tPlqT2t2v+OgvqZhuzI0w5C7Lf
Ap3py/iUoa/RNYfMARaqikdbqiTYMB6G0OoGg4Od/mUkOG5m3fF2BljhrDZnUOnT
04ofmxt5iZLGgBmbPctIUf9iZYMHEi99WYTJpQfHlMYT/ApgQEE8O5YSgNsuNXpO
2g+3aicdmDXeLqJgDMY0JyA6FsnIpNxeKPD0cNdBY32JTQ9daGa4PLbKGMHx8eIe
XsLoUtUDIWF1lTaTq7kgSnmgbelXLI8Db7TcTUoulFNN4MzKLubTuSSG7QaVce2x
fTEVki8xMwvOFoffZQhKLgZZ4A4ya3hhEAKEzg7//dHtmFFI0uq0MQF5pkXZd3JG
osqlSOdLKzbZa/ALM2bRkO4jJZ3ZFF/+9bng2+5WzBZxeYcqgR0yG4bmmGdPyVyf
8axFfeFr2N1X3dyTRtwjRpKknXJbTMT5E5etWAN9tQEX0+fkw/fw0NtBEpVdJAPM
2vRGjYikV0wjNbSOrCw0xjqGImcQD4QX69N+I//aQ5SQfJ0DG9UeVmxFqqnrdaWk
H6GK8/YGfG9k86+eR+0VvBmqzFb+axyxxPRJBlygdwDE6FlLz1xdcuHieStO9Gpz
UUDC8ddo3VxibOWdDXNhodYcGHSwFz9G8QIzxQNubsO5Hw1UR9b+1ba1DjBS07FD
BzVr6f/QsX7MPc1yoftun+UMOaIjBOSIGq9hCklgKfYygNu6koBQI/ZbFIRB3HNb
XP6rH9dN20lwwHujEquawQfTH8B3bCH7zMUrprJDCfpj1c7JOF/uJhQiojQXbFyR
Xubw3yE/+S1ycVpNvQ5NGaoPDk/5d8LFwEdI1r/5Xlx30Ncr/QihEqoiJVdrW2i1
/3YxNdyLmbbdbGFDprBz/dReLRoOiIdOO5wKGl8GBjwQckqu8GcdZ6aTgxS1N1Sv
DwA8a8I9olUECiu4V4xbzV0Tb6bz6dhCDXibV7B4Muqh0tUDwVieahYWQcJukLWO
NiP5XvBv70LBKEDnJzc6IlIz0ZPThRo5RJgbwQv9XuI0E6JeUJXyC/J/S5iHqJod
4t7XQX7bhWf0nfQoIaNSdnbWATyvAn4pHulaheCTnJwA7MKul6rsUcoRGF9XB0ax
eveS6eX1FSWziR6ydS/Oprr1PpM0TXFFN+TAmSVnGWUYl40RWaYdip8N4ghZjCOQ
oemjKPbBQiqImiaUR+00V0W1puFQ1/n5bdTiYOu/687mECuoTCBUJLERLSnQiRJb
crGbAf9l6K/6FJ9EG2rHIzoVaFv4sZW7ei8jXrbwNyU//tfKniGHnTwPaYTV3A/f
bHt4EKSYCGiUKV991fScT+g2IbiMY+SrZWVQ9O+n7yWXPO3ISq8rWXzKVIrxwrdp
VP7104zEVa/bOcdTzYzCQdrupo/eTeld832dXrVj6S2k35Y7g3TLRp5L1tPdM+K0
TFD/pnYEV8vMpDm+2p2dXGRh6MjLfEpsWBt/4+1V4i4XvcPmpH1KOyNx8lQdEGn8
vbtDRkeIaMxw38ZiVaAKHNTqShf1xCN+HFycbWV8YVMrp1Bu2pA2ghOj1IFdvYqz
/g/GVkcwel8prZvCu3MgZC/rkvxe2u78z3QZjVaYDKm+X93u0GTM3D7MrC5e4vhT
QysAtwADDysR63VLlH7+MDg3UvbKiR16UQorcJ4VM3UtJiGickPsffgldSHxLlsi
+dQvDrved1bNgdiNG0UIRfL9+i8zV+NEg80gLJ7cJvsVx6DtklEoGnV+0gIN2bo+
4ACp+fkBbi3H7fm5+Im0JD5AviFqy5/tw0kEGzIpzKVn8S6qVjYRvnt4vzLn34gy
Ov8WhlQOI2RahT3gAK4vvoXk9bDBqvVpBciqjX59zNsc5aeFsDOeHPIiNvzrce7F
TS4GnlE3Xf/belvqfe5Q3aMg4S4Z//aywRoWgQupvr95vOkNv8tMAjos2f9hekHJ
/PmDTFt3NeVrXYiVFtOqYdMqR9o/ZehITjrOt2M0LJW6I9WHyYsE8zp5iIZ6PdjQ
nih1PGxxr/gprDu3HXDKtMT/W4fifopsBLOJok+BAqrrzI1qy1vu0bb+Jj+jaSfX
BVGCUqBisbrcPKPzpzYJA4SSJMFbapig9ZHFbuZeT3fOHH/B59JFNVCXW9c67wkM
DmS+n2SVzn/Bdu55uysv6/a7uaFEkaU1GdI5I15/p+0RoMqVLUljQU0+hYK9rTGu
JApZie5mQyTy3APZbhg+k1DnHJ5F4J8Q1HwrTRYFnZ5KgTxgbtouVBeRpn4oBld4
geB/xemAVwuhYJpO88sEMM/yneixAgenjfeQi3uQXQd0UHSumnuchlvS+mfcHMj3
e/ykx8dsrJHhwyrz7kuTImueg4RpCe1i7j1dMnSET6R5PP/a9i/Xfm1rVt/zH/wT
kuauWhQg+7kXeLUd+JhyKEP7d7HE+ulGp8NF6xUmlcU9LpHXPf1G5pNOnnama2S7
xizPY8drRWk6b8XUFuuaKqFUobH24VOkQQE5MiPapEFiA3KnOeiXxqnN7BnAJeqZ
FsTD17dH0M11PKrI5UNUeb0aUnrf7E77gfgp+WrlJWOtX6vS+ficWy2Yhyz5Rsgt
EEFdwr4AyEmrflF1dF2L5mFZmR3B/hvNXEXfnF54zaY5A0w5ZY5BllaK9pGCDINC
vhCisfrP1RLCczA6tA/Mq+JF6UCsPEV5lRmaPUkSs8LmRWeSRx7D+qd1NOuOJKBW
GV2XhIMOl/wldUSDP/4LjLIC0BbIWR+p2OMpiXQt3clyYpAaATDkyCsvMUSuVIUj
dSg2luIY9ZaXLHN5ycYS018l/C+T0RcqrAXOAlNr7gKnY7qP/MiPiVwefqb2KgwT
yRF6kVae8GstCp2cQwmylixkpLdxXs2epzNHU7n+cAhb5fBfAgBqG7HypdSTcrUr
MltlOjLG9b92w3vOYBZCEkJa8CnttSbWVoFBLdKC9UrN7Z7lakFudHcBxdZq4kUs
5TWGeS8mqyqQ5znp5bdX2OoE7Jjp0f8AMvUzNnt6SatmoEcTQfQ95lkoHmpe5Zzo
6xjSHbzMCZ7sejlMvN6AkN9YvoE9dSZo3I66aytxShxtZppjpdktSFn/D/6v/Oka
PX6pHXGy/3C6rPgy90MuL3/C7b/dRpvEiuIfRfaMXEjec9fW3ZjnDJpnGGI2oAtS
lIKAyaR69f96+VvbQOt8eCMo1q7S9gq70C8OcWe5D+aPj92F3+TXO8IpnrimDCLj
IEikQFV7dUtFQNEulMM5BSRZ34BLwP4dlGP+6m37/dqg+2z5NoVJDw79Bk76L1Yj
8b1kMVZmPDJEGuNklTG17nRNZtf1qyqty/ypLqjUnyJoD1cLTp5DcjcMQPgNLPmZ
Uv8fQaZrDuJZKeldyUfbJAG+k8CE3y0tz4cA+UVDptmXZEHIqhoOnQ0i5pyFbTdA
ShPyi+RJOomyy2M+BcN5MeVumJ/ndiuIB1mi8C7IZR7MNgM0khHrIulXAl9/iR9w
eVJxNbMDKHAJoS47wv5vE+YR32x8UZdL4LMM3jDfYvj4AvrorYQHmrYyQyUPwRNr
bgO8dUHNaz9XKviwbsCMvCgoIT7si+RtnLZeeA+NDJfJRRFuxHPKiLhgeQyUrJav
bBBrr2BkvKMywJCzvxmur+Bwo6Ktl/kc/ZBnq1TXNFLDXxSlY9Uqjf0h7Dbv6/W5
IYmhEjdAocP4HSVgcPM1qFSe8K72mbKzKxtXN0Q3PjDLnys4XbKI5EilvayKHj33
1f/RFMj511+JfkrmaQceSkXAIKK+BPAooi+VvvON5N+uPH6O3LQuvv4ICX00g1lg
LWBKPiQFga3scu/JCci1m8Ao6fBau7n19lmRoysaW/RxlFqn4zsTkiMtNCCmoLMD
jcMCqwM5hISuvSiJXkCM+wgsNpiacZO4c28Y9kYSzA8BGT8lrPLB3GX/5pMlpx1W
6lF2c0TAfe83dWum5OG2oCpqwb04TGzOUVuIk82/S53OrRtEcCiDXxu6d+1oJVDk
edtZ3IF74BWij9P5JUoA2b6+6TrOV3Y4RNlsvjfRg6LmxifS36qu2uERccTgzy74
Jw92hiZKU0n/TXXBb4uJIaJhASxFIcazZCQwZTtekQ6zkVwsvHOX5oRSokuHx03Y
jkcg6Q98Pei1Xh+LYZH7NUR5+nRS4D/32GT2riCG3lBy3xsp3OBJ237q/aPvTTiQ
Uq2ZPUKVU6/QPQLJaAM+T/OO9/it1rSDgJtqFpMXSnPv8VyLzmwO0wwPFUNI8N72
RdGvWh1Tiq9GEnVJ0BcXbiqyK8nCbMVzCJtARxQ7Idwq+MPmDMZnbz5gVZ14SFA7
khpjjTL/TQgnh9sEzdu3Mqmcmj7Ezn8aV8f4CfqzgQZlKlkMBOe+piSkOpHyrD/Q
/fIjJjTbBnWcLAzDjvvgJSwDRF8HlVM8HnLldKVKf2NDvVxBvCxbB+ZXhF9A+wkK
ViY+m6Tt6y8l1cMrWTAq3CX8m6ijgBxwtO+ZWL95IlVTj0tiQFTnT9/4hhJiD2qn
16wfoLiGcJxtBqYGyayEAvqXtAFaZYMO0boeu4BP6yhfuLDBm+WpUe3CODuOjsCF
KrFkW7Y2G6PYQCPL4rTVg2ejI+ETgJpL/vqimX1nvwU3dcyFXJnIqEUgP0djP/Yp
s1i+ItnLFg50uYtmnOsKya5rsznHcT30i4q01qvko9yHq3URaRCE3JkCDeGqojMR
1TR9IeYBoe7EyZnLvqbmHTzzr+r+9n5dqDTBFPNyT+svPmauecBby6XAQgtq//qz
4FsLArxvUIuv0SBtCwGpM+OPWJrwTRucaz9iPWlEz/KocSe00MO0mzyfQuitixPu
e4r2D3RvLlDENmkByQCJqy1EYUvMUIcb+Fu4VNLKA7naeOgwktCvI/xIRSjFLuI6
ZvSYgyC203tEqquAm3RvXgqZDN44ofeYsPxH87f0wTfjuKIm21D1scPqarroE4t+
rvF0u4X3zSfHuGm6yyipEH561VaxMlugogpfwQVvXXz56f4zfU9Mt5V0Ci0Jnzgs
m1b9am51yY74AZQxCPBkXzMH91LJYhUapSSD50/2wkwM0mzrFZJI+7ktqA3mFIyv
st8Vs0A336iubKaHy5Py0eF3DEc6Uvs+1WwzIu4dH1uJ2Y0huKxh/wflGw7wQ4Lq
pS7S2rRVUBXtwEqa2l2+7d2AUl109eK/BqxZF3JX2tCI1ExxD7PLlLcfI2Z8xBNY
RJ9LlOJ7fdgknHdOvrKoFKy0YiQewnjbKE4GRJoXgUyn4hYIjIU5AHkclSYSVHzV
+BjiX/JOZEbVmrSlIoNbNoECt/ndfU31QHsAe0Rx6U+rjPH4IykCWwWQlEb7dKls
TarcBWgMht9GmLdo0bN/BPbOLAD3Y3Utzk+qpKCXJs993r7/cetyto0LQLzRxpxT
JHza4Hk4rhQhNAxusTsSTzA0PcRppwfAGxjb56HQAb2kTj8uZnTj+yXaaRZNWRkj
ocHOMBlB6imugNo1QNVy2lyhw3WUpP25kNGyWz8Km4nsQ7tX6MnRyS+riDwecaI3
/mSvbohQqnjZfTnuYqPP5iN4IRi+B7SkPNrLtHCZfpOOkZLtSrKssbcck+tB2SzI
FgNNyCmpK6eBREbFM5mHPKTSMOj2kc5mM7HLxlzu7TKhjcY/A8ZrUmX3aMfmolEI
kh8tzw1Uxoqg+wFC2aGAK9DJro+9SsiEJ+MBDcvk5xIgU3jhw4BKn0ec0x86UWja
r1P9DF3i4He64Pwn2pYdnIFt6zpsciE+THUSvnwyRd0+seUYH3cjrsS0MC2EDprY
NT9H1a5COBZLiWkjai4bvbBD2NDyLLRzPbQ+8V99MmFbHoDA6QRF/eo6I47JcqAo
fYv9OzmPsccHxRdaNsafmbRqXxLaXJHR0qNrS3nPPh3xpy5Q3axMC8hkmplz17fy
/efRF1Zl5JbsJVE6ccjXgY4HpJTJW9xP0o3MD9V207wy+mOu8rpOgdpisCfYhtWl
SUaWn51ixphdkexpqCLHwNmqfmdXRaE28cn3sYlG1w/1ZZ3I+86sLKN3OIyRqat8
cxrkHwUyiyMFRhcjZ3D0bo2U2e+ZIzxYy3XltzGNVZ9h/VKFsGAVsMs9Ykt7uuyU
xcjISiC96pmfi0f1CLFuEF089jXAI/aPH0mCPm14YsdL5Jdzqc27YeostfAAZ3Hc
GLHJtZLJQ8fE5yrdHhqO6pHKbB9S5dP/8M3OInt2Il3X/an57tqhkCZBNttMKBF9
OhFI4rqlVjpxrKe6/nA/H06oAqxXZXymMOdUfKYBPGZx7mxZKxnoxArUbqBdTAvn
NjXyOAPL1KmFr4QH2AUGrPMEiWlG1P7nUxyE2wRla/zbz5TXZvDCptnf87n56xa1
v3Ne/N0BRFz9mfJb7EfRRc3vbEqjNSO0V4x4zbciHF0y/bkQ9v5Odmyq6Nk6Aoxn
altn+XxKDAJGWPj8JXqOWrGTH1xhM9N04yz9R80giR0Mekrs/fy6NGqzrIiVU0Jb
wfLF1UP2ILnY9Kzh/6IBW121jvYvFp6LaQLGlcO1XDUFL1Aogm6xyED3VjMeMPVs
90dYDN669e4IpJi43vaEcKiQkVoFhGMeBiOrVPsvNKmqGdgLhvkP7fwEGQPmG9St
I0nzaxZElkK2or5C+SS9gML2NTw00BfEP+o272cx0ZiXSElqgUVIDF41lD75tNvU
lCekwkpkqgG1P+Wgt4IMsXwqnSEJlsH1NY7jpozFY7UIn1vRubyY/J9PU4APGC4E
ya5jP9bL6abhE1caDL43H44rP/0FGC/wtwcvQm7cXrbfB50Vv7eo8Oe8gYmp26wI
LOmfvxzcORrekbgr3OQxtdrvzz0x+DEhBap5x6cbBZZmLD33T18fDbYzgcpBU84W
owQ9b0pHHK/w65c9Q9oNZvLm9Y6X8GRryM75P2WI0e/0aRfXYoitXcXBiAxf1BoV
UZK53o12Utxwu7Iva459Cru2knhH4RDohGeMpAGMErBL8378NOrR0ZEUHL/vh1ab
Y6AJEvqeJHQiBB3QGJjfLglnfQvK0HGBZfBpvecuZNa/OcXGyd4ubD9oNQbBaB+1
6Dn1/yoCzWI5d2sqtKOJHMRiUuknAsLGjLMxlGjfyhdn5ydOJsYTJ4Oz8kAXygMm
t5z0NrZ/jwjUvmZl++2136QGMgBdHOQ99cUAT3l6k6VDU7oPcZ6l0xp58w1IwxaN
OeZFZyZwPbW5nf5hploD9Qua8NtKlB7yBgQh81zjAOWkmO/2NKO6XyqMqziIqZRq
iDi8QzBkg1SqKF7RwuUxMaZittBf5GKf12BNRX0A913z+iLDTim7xaV+i6nzGVXv
4jHoCBG0rT5L+5l3hpFmzJ4/qOf360twUE4VtDePLoD9JSqlNgumVtWgOQGYpF1l
j6tCnlfIquHttKPipVNw9okorBFdmc00akcI1XyCNomcn4gIsTfoT71aGo2HjTPJ
FO4CviW9axp3yjKwEj5kczkghBi29xw0GIHLTIuAHNP8nSeQI1GfNchBTgNYD8di
Ceexwq89u+b01K1RL4LJJc/HWD9FPv9B8E/mqd4OzdiuguVZ0x5sz2GA5sIXBgvs
ZjSoh3myVbIbIHx3xOJN86y8estLTZzGvivItyzIH067mzlzpqicRWIqF5+gQdVE
vQcZh+qG3ZXLddg6P/FsFPxr+W/wQUEMzwJ4AJVL8Fo=
`pragma protect end_protected
